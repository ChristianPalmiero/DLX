
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_dataPath is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_dataPath;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Adder_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Adder_DW01_add_0;

architecture SYN_rpl of Adder_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, net88777 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           net88777, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity comparator_DW01_cmp6_1 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_DW01_cmp6_1;

architecture SYN_rpl of comparator_DW01_cmp6_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47 : std_logic;

begin
   
   U19 : XOR2_X1 port map( A => B(10), B => A(10), Z => n23);
   U20 : XOR2_X1 port map( A => B(9), B => A(9), Z => n22);
   U21 : XOR2_X1 port map( A => B(8), B => A(8), Z => n21);
   U22 : XOR2_X1 port map( A => B(7), B => A(7), Z => n20);
   U24 : XOR2_X1 port map( A => B(14), B => A(14), Z => n27);
   U25 : XOR2_X1 port map( A => B(13), B => A(13), Z => n26);
   U26 : XOR2_X1 port map( A => B(12), B => A(12), Z => n25);
   U27 : XOR2_X1 port map( A => B(11), B => A(11), Z => n24);
   U30 : XOR2_X1 port map( A => B(18), B => A(18), Z => n35);
   U31 : XOR2_X1 port map( A => B(17), B => A(17), Z => n34);
   U32 : XOR2_X1 port map( A => B(16), B => A(16), Z => n33);
   U33 : XOR2_X1 port map( A => B(15), B => A(15), Z => n32);
   U35 : XOR2_X1 port map( A => B(22), B => A(22), Z => n39);
   U36 : XOR2_X1 port map( A => B(21), B => A(21), Z => n38);
   U37 : XOR2_X1 port map( A => B(20), B => A(20), Z => n37);
   U38 : XOR2_X1 port map( A => B(19), B => A(19), Z => n36);
   U40 : XOR2_X1 port map( A => B(26), B => A(26), Z => n43);
   U41 : XOR2_X1 port map( A => B(25), B => A(25), Z => n42);
   U42 : XOR2_X1 port map( A => B(24), B => A(24), Z => n41);
   U43 : XOR2_X1 port map( A => B(23), B => A(23), Z => n40);
   U45 : XOR2_X1 port map( A => B(30), B => A(30), Z => n47);
   U46 : XOR2_X1 port map( A => B(29), B => A(29), Z => n46);
   U47 : XOR2_X1 port map( A => B(28), B => A(28), Z => n45);
   U48 : XOR2_X1 port map( A => B(27), B => A(27), Z => n44);
   U1 : NOR4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => EQ);
   U2 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n2);
   U3 : NAND4_X1 port map( A1 => n5, A2 => n6, A3 => n7, A4 => n8, ZN => n4);
   U4 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => n1
                           );
   U5 : NOR4_X1 port map( A1 => n44, A2 => n45, A3 => n46, A4 => n47, ZN => n28
                           );
   U6 : NOR4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => n29
                           );
   U7 : NOR4_X1 port map( A1 => n36, A2 => n37, A3 => n38, A4 => n39, ZN => n30
                           );
   U8 : NOR4_X1 port map( A1 => n32, A2 => n33, A3 => n34, A4 => n35, ZN => n31
                           );
   U9 : NOR4_X1 port map( A1 => n20, A2 => n21, A3 => n22, A4 => n23, ZN => n19
                           );
   U10 : NOR4_X1 port map( A1 => n24, A2 => n25, A3 => n26, A4 => n27, ZN => 
                           n18);
   U11 : OAI22_X1 port map( A1 => n13, A2 => n14, B1 => B(1), B2 => n13, ZN => 
                           n12);
   U12 : INV_X1 port map( A => A(1), ZN => n14);
   U13 : AND2_X1 port map( A1 => B(0), A2 => n15, ZN => n13);
   U14 : NOR2_X1 port map( A1 => n15, A2 => B(0), ZN => n16);
   U15 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n8);
   U16 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n7);
   U17 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n6);
   U18 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n3
                           );
   U23 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n9);
   U28 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n10);
   U29 : OAI22_X1 port map( A1 => A(1), A2 => n16, B1 => n16, B2 => n17, ZN => 
                           n11);
   U34 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n5);
   U39 : INV_X1 port map( A => A(0), ZN => n15);
   U44 : INV_X1 port map( A => B(1), ZN => n17);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity comparator_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end comparator_DW01_cmp6_0;

architecture SYN_rpl of comparator_DW01_cmp6_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n201, n202, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200 : std_logic;

begin
   
   U24 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => n68);
   U25 : NAND3_X1 port map( A1 => n74, A2 => n75, A3 => n76, ZN => n71);
   U42 : XOR2_X1 port map( A => n99, B => B(30), Z => n7);
   U1 : INV_X1 port map( A => n59, ZN => n167);
   U2 : INV_X1 port map( A => n39, ZN => n139);
   U3 : INV_X1 port map( A => n19, ZN => n111);
   U4 : AOI211_X1 port map( C1 => n67, C2 => n68, A => n69, B => n70, ZN => n61
                           );
   U5 : NOR2_X1 port map( A1 => n83, A2 => n84, ZN => n67);
   U6 : AOI211_X1 port map( C1 => n57, C2 => n58, A => n59, B => n60, ZN => n51
                           );
   U7 : NOR2_X1 port map( A1 => n85, A2 => n86, ZN => n57);
   U8 : OAI211_X1 port map( C1 => n61, C2 => n62, A => n63, B => n64, ZN => n58
                           );
   U9 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => n62);
   U10 : AOI211_X1 port map( C1 => n47, C2 => n48, A => n49, B => n50, ZN => 
                           n41);
   U11 : NOR2_X1 port map( A1 => n87, A2 => n88, ZN => n47);
   U12 : OAI211_X1 port map( C1 => n51, C2 => n52, A => n53, B => n54, ZN => 
                           n48);
   U13 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => n52);
   U14 : AOI211_X1 port map( C1 => n37, C2 => n38, A => n39, B => n40, ZN => 
                           n31);
   U15 : NOR2_X1 port map( A1 => n89, A2 => n90, ZN => n37);
   U16 : OAI211_X1 port map( C1 => n41, C2 => n42, A => n43, B => n44, ZN => 
                           n38);
   U17 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => n42);
   U18 : AOI211_X1 port map( C1 => n27, C2 => n28, A => n29, B => n30, ZN => 
                           n21);
   U19 : NOR2_X1 port map( A1 => n91, A2 => n92, ZN => n27);
   U20 : OAI211_X1 port map( C1 => n31, C2 => n32, A => n33, B => n34, ZN => 
                           n28);
   U21 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => n32);
   U22 : AOI211_X1 port map( C1 => n17, C2 => n18, A => n19, B => n20, ZN => 
                           n11);
   U23 : NOR2_X1 port map( A1 => n93, A2 => n94, ZN => n17);
   U26 : OAI211_X1 port map( C1 => n21, C2 => n22, A => n23, B => n24, ZN => 
                           n18);
   U27 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n22);
   U28 : NOR2_X1 port map( A1 => n195, A2 => n196, ZN => n79);
   U29 : INV_X1 port map( A => n75, ZN => n196);
   U30 : NOR2_X1 port map( A1 => n175, A2 => n85, ZN => n64);
   U31 : NOR2_X1 port map( A1 => n161, A2 => n87, ZN => n54);
   U32 : NOR2_X1 port map( A1 => n147, A2 => n89, ZN => n44);
   U33 : NOR2_X1 port map( A1 => n133, A2 => n91, ZN => n34);
   U34 : NOR2_X1 port map( A1 => n119, A2 => n93, ZN => n24);
   U35 : NOR2_X1 port map( A1 => n105, A2 => n95, ZN => n14);
   U36 : AOI21_X1 port map( B1 => n171, B2 => n172, A => n86, ZN => n166);
   U37 : INV_X1 port map( A => n60, ZN => n172);
   U38 : AOI21_X1 port map( B1 => n174, B2 => n64, A => n175, ZN => n171);
   U39 : AOI21_X1 port map( B1 => n177, B2 => n63, A => n178, ZN => n174);
   U40 : AOI21_X1 port map( B1 => n143, B2 => n144, A => n90, ZN => n138);
   U41 : INV_X1 port map( A => n40, ZN => n144);
   U43 : AOI21_X1 port map( B1 => n146, B2 => n44, A => n147, ZN => n143);
   U44 : AOI21_X1 port map( B1 => n149, B2 => n43, A => n150, ZN => n146);
   U45 : AOI21_X1 port map( B1 => n115, B2 => n116, A => n94, ZN => n110);
   U46 : INV_X1 port map( A => n20, ZN => n116);
   U47 : AOI21_X1 port map( B1 => n118, B2 => n24, A => n119, ZN => n115);
   U48 : AOI21_X1 port map( B1 => n121, B2 => n23, A => n122, ZN => n118);
   U49 : AOI21_X1 port map( B1 => n188, B2 => n73, A => n189, ZN => n185);
   U50 : AOI21_X1 port map( B1 => n191, B2 => n72, A => n192, ZN => n188);
   U51 : INV_X1 port map( A => n74, ZN => n192);
   U52 : AOI21_X1 port map( B1 => n194, B2 => n79, A => n195, ZN => n191);
   U53 : AOI21_X1 port map( B1 => n180, B2 => n181, A => n182, ZN => n177);
   U54 : INV_X1 port map( A => n69, ZN => n181);
   U55 : AOI21_X1 port map( B1 => n185, B2 => n186, A => n84, ZN => n180);
   U56 : INV_X1 port map( A => n70, ZN => n186);
   U57 : AOI21_X1 port map( B1 => n160, B2 => n54, A => n161, ZN => n157);
   U58 : AOI21_X1 port map( B1 => n163, B2 => n53, A => n164, ZN => n160);
   U59 : INV_X1 port map( A => n55, ZN => n164);
   U60 : AOI21_X1 port map( B1 => n166, B2 => n167, A => n168, ZN => n163);
   U61 : AOI21_X1 port map( B1 => n152, B2 => n153, A => n154, ZN => n149);
   U62 : INV_X1 port map( A => n49, ZN => n153);
   U63 : AOI21_X1 port map( B1 => n157, B2 => n158, A => n88, ZN => n152);
   U64 : INV_X1 port map( A => n50, ZN => n158);
   U65 : AOI21_X1 port map( B1 => n132, B2 => n34, A => n133, ZN => n129);
   U66 : AOI21_X1 port map( B1 => n135, B2 => n33, A => n136, ZN => n132);
   U67 : INV_X1 port map( A => n35, ZN => n136);
   U68 : AOI21_X1 port map( B1 => n138, B2 => n139, A => n140, ZN => n135);
   U69 : AOI21_X1 port map( B1 => n124, B2 => n125, A => n126, ZN => n121);
   U70 : INV_X1 port map( A => n29, ZN => n125);
   U71 : AOI21_X1 port map( B1 => n129, B2 => n130, A => n92, ZN => n124);
   U72 : INV_X1 port map( A => n30, ZN => n130);
   U73 : AOI21_X1 port map( B1 => n104, B2 => n14, A => n105, ZN => n101);
   U74 : AOI21_X1 port map( B1 => n107, B2 => n13, A => n108, ZN => n104);
   U75 : INV_X1 port map( A => n15, ZN => n108);
   U76 : AOI21_X1 port map( B1 => n110, B2 => n111, A => n112, ZN => n107);
   U77 : AOI21_X1 port map( B1 => n8, B2 => n9, A => n10, ZN => n6);
   U78 : NOR2_X1 port map( A1 => n95, A2 => n96, ZN => n8);
   U79 : OAI211_X1 port map( C1 => n11, C2 => n12, A => n13, B => n14, ZN => n9
                           );
   U80 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => n12);
   U81 : NOR2_X1 port map( A1 => n189, A2 => n83, ZN => n73);
   U82 : NAND2_X1 port map( A1 => n183, A2 => n66, ZN => n69);
   U83 : INV_X1 port map( A => n182, ZN => n183);
   U84 : NAND2_X1 port map( A1 => n169, A2 => n56, ZN => n59);
   U85 : INV_X1 port map( A => n168, ZN => n169);
   U86 : NAND2_X1 port map( A1 => n155, A2 => n46, ZN => n49);
   U87 : INV_X1 port map( A => n154, ZN => n155);
   U88 : NAND2_X1 port map( A1 => n141, A2 => n36, ZN => n39);
   U89 : INV_X1 port map( A => n140, ZN => n141);
   U90 : NAND2_X1 port map( A1 => n127, A2 => n26, ZN => n29);
   U91 : INV_X1 port map( A => n126, ZN => n127);
   U92 : NAND2_X1 port map( A1 => n113, A2 => n16, ZN => n19);
   U93 : INV_X1 port map( A => n112, ZN => n113);
   U94 : INV_X1 port map( A => n10, ZN => n102);
   U95 : INV_X1 port map( A => n65, ZN => n178);
   U96 : INV_X1 port map( A => n45, ZN => n150);
   U97 : INV_X1 port map( A => n25, ZN => n122);
   U98 : NOR2_X1 port map( A1 => n187, A2 => A(5), ZN => n70);
   U99 : NOR2_X1 port map( A1 => n173, A2 => A(9), ZN => n60);
   U100 : NOR2_X1 port map( A1 => n159, A2 => A(13), ZN => n50);
   U101 : NOR2_X1 port map( A1 => n145, A2 => A(17), ZN => n40);
   U102 : NOR2_X1 port map( A1 => n131, A2 => A(21), ZN => n30);
   U103 : NOR2_X1 port map( A1 => n117, A2 => A(25), ZN => n20);
   U104 : NOR2_X1 port map( A1 => n197, A2 => A(2), ZN => n195);
   U105 : NOR2_X1 port map( A1 => n190, A2 => A(4), ZN => n189);
   U106 : NOR2_X1 port map( A1 => n176, A2 => A(8), ZN => n175);
   U107 : NOR2_X1 port map( A1 => n162, A2 => A(12), ZN => n161);
   U108 : NOR2_X1 port map( A1 => n148, A2 => A(16), ZN => n147);
   U109 : NOR2_X1 port map( A1 => n134, A2 => A(20), ZN => n133);
   U110 : NOR2_X1 port map( A1 => n120, A2 => A(24), ZN => n119);
   U111 : NOR2_X1 port map( A1 => n106, A2 => A(28), ZN => n105);
   U112 : NOR2_X1 port map( A1 => n184, A2 => A(6), ZN => n182);
   U113 : NOR2_X1 port map( A1 => n170, A2 => A(10), ZN => n168);
   U114 : NOR2_X1 port map( A1 => n156, A2 => A(14), ZN => n154);
   U115 : NOR2_X1 port map( A1 => n142, A2 => A(18), ZN => n140);
   U116 : NOR2_X1 port map( A1 => n128, A2 => A(22), ZN => n126);
   U117 : NOR2_X1 port map( A1 => n114, A2 => A(26), ZN => n112);
   U118 : NOR2_X1 port map( A1 => n103, A2 => A(29), ZN => n10);
   U119 : NOR2_X1 port map( A1 => n98, A2 => A(31), ZN => n3);
   U120 : OAI211_X1 port map( C1 => A(1), C2 => n77, A => n78, B => n79, ZN => 
                           n76);
   U121 : INV_X1 port map( A => n81, ZN => n77);
   U122 : OAI21_X1 port map( B1 => n80, B2 => n81, A => B(1), ZN => n78);
   U123 : NAND2_X1 port map( A1 => A(0), A2 => n82, ZN => n81);
   U124 : NAND2_X1 port map( A1 => A(6), A2 => n184, ZN => n66);
   U125 : NAND2_X1 port map( A1 => A(10), A2 => n170, ZN => n56);
   U126 : NAND2_X1 port map( A1 => A(14), A2 => n156, ZN => n46);
   U127 : NAND2_X1 port map( A1 => A(18), A2 => n142, ZN => n36);
   U128 : NAND2_X1 port map( A1 => A(22), A2 => n128, ZN => n26);
   U129 : NAND2_X1 port map( A1 => A(26), A2 => n114, ZN => n16);
   U130 : NAND2_X1 port map( A1 => A(31), A2 => n98, ZN => n1);
   U131 : NAND2_X1 port map( A1 => A(7), A2 => n179, ZN => n65);
   U132 : NAND2_X1 port map( A1 => A(11), A2 => n165, ZN => n55);
   U133 : NAND2_X1 port map( A1 => A(15), A2 => n151, ZN => n45);
   U134 : NAND2_X1 port map( A1 => A(19), A2 => n137, ZN => n35);
   U135 : NAND2_X1 port map( A1 => A(23), A2 => n123, ZN => n25);
   U136 : NAND2_X1 port map( A1 => A(27), A2 => n109, ZN => n15);
   U137 : INV_X1 port map( A => A(1), ZN => n80);
   U138 : AND2_X1 port map( A1 => A(4), A2 => n190, ZN => n83);
   U139 : AND2_X1 port map( A1 => A(8), A2 => n176, ZN => n85);
   U140 : AND2_X1 port map( A1 => A(12), A2 => n162, ZN => n87);
   U141 : AND2_X1 port map( A1 => A(16), A2 => n148, ZN => n89);
   U142 : AND2_X1 port map( A1 => A(20), A2 => n134, ZN => n91);
   U143 : AND2_X1 port map( A1 => A(24), A2 => n120, ZN => n93);
   U144 : AND2_X1 port map( A1 => A(28), A2 => n106, ZN => n95);
   U145 : AND2_X1 port map( A1 => A(5), A2 => n187, ZN => n84);
   U146 : AND2_X1 port map( A1 => A(9), A2 => n173, ZN => n86);
   U147 : AND2_X1 port map( A1 => A(13), A2 => n159, ZN => n88);
   U148 : AND2_X1 port map( A1 => A(17), A2 => n145, ZN => n90);
   U149 : AND2_X1 port map( A1 => A(21), A2 => n131, ZN => n92);
   U150 : AND2_X1 port map( A1 => A(25), A2 => n117, ZN => n94);
   U151 : AND2_X1 port map( A1 => A(29), A2 => n103, ZN => n96);
   U152 : OR2_X1 port map( A1 => n179, A2 => A(7), ZN => n63);
   U153 : OR2_X1 port map( A1 => n165, A2 => A(11), ZN => n53);
   U154 : OR2_X1 port map( A1 => n151, A2 => A(15), ZN => n43);
   U155 : OR2_X1 port map( A1 => n137, A2 => A(19), ZN => n33);
   U156 : OR2_X1 port map( A1 => n123, A2 => A(23), ZN => n23);
   U157 : OR2_X1 port map( A1 => n109, A2 => A(27), ZN => n13);
   U158 : NAND2_X1 port map( A1 => A(2), A2 => n197, ZN => n75);
   U159 : NAND2_X1 port map( A1 => A(3), A2 => n193, ZN => n74);
   U160 : INV_X1 port map( A => n201, ZN => GE);
   U161 : OAI21_X1 port map( B1 => n3, B2 => n97, A => n1, ZN => n201);
   U162 : AOI22_X1 port map( A1 => B(30), A2 => n99, B1 => n100, B2 => n7, ZN 
                           => n97);
   U163 : AOI21_X1 port map( B1 => n101, B2 => n102, A => n96, ZN => n100);
   U164 : INV_X1 port map( A => n202, ZN => GT);
   U165 : AOI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => n202);
   U166 : INV_X1 port map( A => n4, ZN => n2);
   U167 : AOI22_X1 port map( A1 => A(30), A2 => n5, B1 => n6, B2 => n7, ZN => 
                           n4);
   U168 : INV_X1 port map( A => B(2), ZN => n197);
   U169 : INV_X1 port map( A => B(6), ZN => n184);
   U170 : INV_X1 port map( A => B(10), ZN => n170);
   U171 : INV_X1 port map( A => B(14), ZN => n156);
   U172 : INV_X1 port map( A => B(0), ZN => n82);
   U173 : INV_X1 port map( A => B(18), ZN => n142);
   U174 : INV_X1 port map( A => B(22), ZN => n128);
   U175 : INV_X1 port map( A => B(26), ZN => n114);
   U176 : INV_X1 port map( A => B(31), ZN => n98);
   U177 : OR2_X1 port map( A1 => n193, A2 => A(3), ZN => n72);
   U178 : INV_X1 port map( A => A(30), ZN => n99);
   U179 : INV_X1 port map( A => B(3), ZN => n193);
   U180 : INV_X1 port map( A => B(7), ZN => n179);
   U181 : INV_X1 port map( A => B(11), ZN => n165);
   U182 : INV_X1 port map( A => B(15), ZN => n151);
   U183 : INV_X1 port map( A => B(19), ZN => n137);
   U184 : INV_X1 port map( A => B(23), ZN => n123);
   U185 : INV_X1 port map( A => B(27), ZN => n109);
   U186 : INV_X1 port map( A => B(4), ZN => n190);
   U187 : INV_X1 port map( A => B(5), ZN => n187);
   U188 : INV_X1 port map( A => B(8), ZN => n176);
   U189 : INV_X1 port map( A => B(9), ZN => n173);
   U190 : INV_X1 port map( A => B(12), ZN => n162);
   U191 : INV_X1 port map( A => B(13), ZN => n159);
   U192 : INV_X1 port map( A => B(16), ZN => n148);
   U193 : INV_X1 port map( A => B(17), ZN => n145);
   U194 : INV_X1 port map( A => B(20), ZN => n134);
   U195 : INV_X1 port map( A => B(21), ZN => n131);
   U196 : INV_X1 port map( A => B(25), ZN => n117);
   U197 : INV_X1 port map( A => B(24), ZN => n120);
   U198 : INV_X1 port map( A => B(28), ZN => n106);
   U199 : INV_X1 port map( A => B(29), ZN => n103);
   U200 : INV_X1 port map( A => n198, ZN => n194);
   U201 : OAI22_X1 port map( A1 => n199, A2 => B(1), B1 => n80, B2 => n200, ZN 
                           => n198);
   U202 : AND2_X1 port map( A1 => n200, A2 => n80, ZN => n199);
   U203 : NOR2_X1 port map( A1 => n82, A2 => A(0), ZN => n200);
   U204 : INV_X1 port map( A => B(30), ZN => n5);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Shifter_NBIT32_DW_rbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_NBIT32_DW_rbsh_0;

architecture SYN_mx2 of Shifter_NBIT32_DW_rbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal MR_int_1_31_port, MR_int_1_30_port, MR_int_1_29_port, 
      MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, MR_int_1_25_port, 
      MR_int_1_24_port, MR_int_1_23_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_20_port, MR_int_1_19_port, MR_int_1_18_port, MR_int_1_17_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_1_0_port, MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, 
      MR_int_2_28_port, MR_int_2_27_port, MR_int_2_26_port, MR_int_2_25_port, 
      MR_int_2_24_port, MR_int_2_23_port, MR_int_2_22_port, MR_int_2_21_port, 
      MR_int_2_20_port, MR_int_2_19_port, MR_int_2_18_port, MR_int_2_17_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_14_port, MR_int_2_13_port, 
      MR_int_2_12_port, MR_int_2_11_port, MR_int_2_10_port, MR_int_2_9_port, 
      MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, MR_int_2_5_port, 
      MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, MR_int_2_1_port, 
      MR_int_2_0_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_28_port, MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, 
      MR_int_3_24_port, MR_int_3_23_port, MR_int_3_22_port, MR_int_3_21_port, 
      MR_int_3_20_port, MR_int_3_19_port, MR_int_3_18_port, MR_int_3_17_port, 
      MR_int_3_16_port, MR_int_3_15_port, MR_int_3_14_port, MR_int_3_13_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_5_port, 
      MR_int_3_4_port, MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, 
      MR_int_3_0_port, MR_int_4_31_port, MR_int_4_30_port, MR_int_4_29_port, 
      MR_int_4_28_port, MR_int_4_27_port, MR_int_4_26_port, MR_int_4_25_port, 
      MR_int_4_24_port, MR_int_4_23_port, MR_int_4_22_port, MR_int_4_21_port, 
      MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, MR_int_4_17_port, 
      MR_int_4_16_port, MR_int_4_15_port, MR_int_4_14_port, MR_int_4_13_port, 
      MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, MR_int_4_9_port, 
      MR_int_4_8_port, MR_int_4_7_port, MR_int_4_6_port, MR_int_4_5_port, 
      MR_int_4_4_port, MR_int_4_3_port, MR_int_4_2_port, MR_int_4_1_port, 
      MR_int_4_0_port, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => MR_int_4_31_port, B => MR_int_4_15_port, S 
                           => n42, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => MR_int_4_30_port, B => MR_int_4_14_port, S 
                           => n42, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => MR_int_4_29_port, B => MR_int_4_13_port, S 
                           => n42, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => MR_int_4_28_port, B => MR_int_4_12_port, S 
                           => n42, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => MR_int_4_27_port, B => MR_int_4_11_port, S 
                           => n42, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => MR_int_4_26_port, B => MR_int_4_10_port, S 
                           => n42, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => MR_int_4_25_port, B => MR_int_4_9_port, S 
                           => n42, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => MR_int_4_24_port, B => MR_int_4_8_port, S 
                           => n42, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => MR_int_4_23_port, B => MR_int_4_7_port, S 
                           => n41, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => MR_int_4_22_port, B => MR_int_4_6_port, S 
                           => n41, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => MR_int_4_21_port, B => MR_int_4_5_port, S 
                           => n41, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => MR_int_4_20_port, B => MR_int_4_4_port, S 
                           => n41, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => MR_int_4_19_port, B => MR_int_4_3_port, S 
                           => n41, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => MR_int_4_18_port, B => MR_int_4_2_port, S 
                           => n41, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => MR_int_4_17_port, B => MR_int_4_1_port, S 
                           => n41, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => MR_int_4_16_port, B => MR_int_4_0_port, S 
                           => n41, Z => B(16));
   M1_4_15 : MUX2_X1 port map( A => MR_int_4_15_port, B => MR_int_4_31_port, S 
                           => n41, Z => B(15));
   M1_4_14 : MUX2_X1 port map( A => MR_int_4_14_port, B => MR_int_4_30_port, S 
                           => n41, Z => B(14));
   M1_4_13 : MUX2_X1 port map( A => MR_int_4_13_port, B => MR_int_4_29_port, S 
                           => n41, Z => B(13));
   M1_4_12 : MUX2_X1 port map( A => MR_int_4_12_port, B => MR_int_4_28_port, S 
                           => n41, Z => B(12));
   M1_4_11 : MUX2_X1 port map( A => MR_int_4_11_port, B => MR_int_4_27_port, S 
                           => n40, Z => B(11));
   M1_4_10 : MUX2_X1 port map( A => MR_int_4_10_port, B => MR_int_4_26_port, S 
                           => n40, Z => B(10));
   M1_4_9 : MUX2_X1 port map( A => MR_int_4_9_port, B => MR_int_4_25_port, S =>
                           n40, Z => B(9));
   M1_4_8 : MUX2_X1 port map( A => MR_int_4_8_port, B => MR_int_4_24_port, S =>
                           n40, Z => B(8));
   M1_4_7 : MUX2_X1 port map( A => MR_int_4_7_port, B => MR_int_4_23_port, S =>
                           n40, Z => B(7));
   M1_4_6 : MUX2_X1 port map( A => MR_int_4_6_port, B => MR_int_4_22_port, S =>
                           n40, Z => B(6));
   M1_4_5 : MUX2_X1 port map( A => MR_int_4_5_port, B => MR_int_4_21_port, S =>
                           n40, Z => B(5));
   M1_4_4 : MUX2_X1 port map( A => MR_int_4_4_port, B => MR_int_4_20_port, S =>
                           n40, Z => B(4));
   M1_4_3 : MUX2_X1 port map( A => MR_int_4_3_port, B => MR_int_4_19_port, S =>
                           n40, Z => B(3));
   M1_4_2 : MUX2_X1 port map( A => MR_int_4_2_port, B => MR_int_4_18_port, S =>
                           n40, Z => B(2));
   M1_4_1 : MUX2_X1 port map( A => MR_int_4_1_port, B => MR_int_4_17_port, S =>
                           n40, Z => B(1));
   M1_4_0 : MUX2_X1 port map( A => MR_int_4_0_port, B => MR_int_4_16_port, S =>
                           n40, Z => B(0));
   M1_3_31_0 : MUX2_X1 port map( A => MR_int_3_31_port, B => MR_int_3_7_port, S
                           => n39, Z => MR_int_4_31_port);
   M1_3_30_0 : MUX2_X1 port map( A => MR_int_3_30_port, B => MR_int_3_6_port, S
                           => n39, Z => MR_int_4_30_port);
   M1_3_29_0 : MUX2_X1 port map( A => MR_int_3_29_port, B => MR_int_3_5_port, S
                           => n39, Z => MR_int_4_29_port);
   M1_3_28_0 : MUX2_X1 port map( A => MR_int_3_28_port, B => MR_int_3_4_port, S
                           => n39, Z => MR_int_4_28_port);
   M1_3_27_0 : MUX2_X1 port map( A => MR_int_3_27_port, B => MR_int_3_3_port, S
                           => n39, Z => MR_int_4_27_port);
   M1_3_26_0 : MUX2_X1 port map( A => MR_int_3_26_port, B => MR_int_3_2_port, S
                           => n39, Z => MR_int_4_26_port);
   M1_3_25_0 : MUX2_X1 port map( A => MR_int_3_25_port, B => MR_int_3_1_port, S
                           => n39, Z => MR_int_4_25_port);
   M1_3_24_0 : MUX2_X1 port map( A => MR_int_3_24_port, B => MR_int_3_0_port, S
                           => n39, Z => MR_int_4_24_port);
   M1_3_23_0 : MUX2_X1 port map( A => MR_int_3_23_port, B => MR_int_3_31_port, 
                           S => n38, Z => MR_int_4_23_port);
   M1_3_22_0 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, 
                           S => n38, Z => MR_int_4_22_port);
   M1_3_21_0 : MUX2_X1 port map( A => MR_int_3_21_port, B => MR_int_3_29_port, 
                           S => n38, Z => MR_int_4_21_port);
   M1_3_20_0 : MUX2_X1 port map( A => MR_int_3_20_port, B => MR_int_3_28_port, 
                           S => n38, Z => MR_int_4_20_port);
   M1_3_19_0 : MUX2_X1 port map( A => MR_int_3_19_port, B => MR_int_3_27_port, 
                           S => n38, Z => MR_int_4_19_port);
   M1_3_18_0 : MUX2_X1 port map( A => MR_int_3_18_port, B => MR_int_3_26_port, 
                           S => n38, Z => MR_int_4_18_port);
   M1_3_17_0 : MUX2_X1 port map( A => MR_int_3_17_port, B => MR_int_3_25_port, 
                           S => n38, Z => MR_int_4_17_port);
   M1_3_16_0 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_24_port, 
                           S => n38, Z => MR_int_4_16_port);
   M1_3_15_0 : MUX2_X1 port map( A => MR_int_3_15_port, B => MR_int_3_23_port, 
                           S => n38, Z => MR_int_4_15_port);
   M1_3_14_0 : MUX2_X1 port map( A => MR_int_3_14_port, B => MR_int_3_22_port, 
                           S => n38, Z => MR_int_4_14_port);
   M1_3_13_0 : MUX2_X1 port map( A => MR_int_3_13_port, B => MR_int_3_21_port, 
                           S => n38, Z => MR_int_4_13_port);
   M1_3_12_0 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, 
                           S => n38, Z => MR_int_4_12_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => n37, Z => MR_int_4_11_port);
   M1_3_10_0 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, 
                           S => n37, Z => MR_int_4_10_port);
   M1_3_9_0 : MUX2_X1 port map( A => MR_int_3_9_port, B => MR_int_3_17_port, S 
                           => n37, Z => MR_int_4_9_port);
   M1_3_8_0 : MUX2_X1 port map( A => MR_int_3_8_port, B => MR_int_3_16_port, S 
                           => n37, Z => MR_int_4_8_port);
   M1_3_7 : MUX2_X1 port map( A => MR_int_3_7_port, B => MR_int_3_15_port, S =>
                           n37, Z => MR_int_4_7_port);
   M1_3_6 : MUX2_X1 port map( A => MR_int_3_6_port, B => MR_int_3_14_port, S =>
                           n37, Z => MR_int_4_6_port);
   M1_3_5 : MUX2_X1 port map( A => MR_int_3_5_port, B => MR_int_3_13_port, S =>
                           n37, Z => MR_int_4_5_port);
   M1_3_4 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S =>
                           n37, Z => MR_int_4_4_port);
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           n37, Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           n37, Z => MR_int_4_2_port);
   M1_3_1 : MUX2_X1 port map( A => MR_int_3_1_port, B => MR_int_3_9_port, S => 
                           n37, Z => MR_int_4_1_port);
   M1_3_0 : MUX2_X1 port map( A => MR_int_3_0_port, B => MR_int_3_8_port, S => 
                           n37, Z => MR_int_4_0_port);
   M1_2_31_0 : MUX2_X1 port map( A => MR_int_2_31_port, B => MR_int_2_3_port, S
                           => n36, Z => MR_int_3_31_port);
   M1_2_30_0 : MUX2_X1 port map( A => MR_int_2_30_port, B => MR_int_2_2_port, S
                           => n36, Z => MR_int_3_30_port);
   M1_2_29_0 : MUX2_X1 port map( A => MR_int_2_29_port, B => MR_int_2_1_port, S
                           => n36, Z => MR_int_3_29_port);
   M1_2_28_0 : MUX2_X1 port map( A => MR_int_2_28_port, B => MR_int_2_0_port, S
                           => n36, Z => MR_int_3_28_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => n36, Z => MR_int_3_27_port);
   M1_2_26_0 : MUX2_X1 port map( A => MR_int_2_26_port, B => MR_int_2_30_port, 
                           S => n36, Z => MR_int_3_26_port);
   M1_2_25_0 : MUX2_X1 port map( A => MR_int_2_25_port, B => MR_int_2_29_port, 
                           S => n36, Z => MR_int_3_25_port);
   M1_2_24_0 : MUX2_X1 port map( A => MR_int_2_24_port, B => MR_int_2_28_port, 
                           S => n36, Z => MR_int_3_24_port);
   M1_2_23_0 : MUX2_X1 port map( A => MR_int_2_23_port, B => MR_int_2_27_port, 
                           S => n35, Z => MR_int_3_23_port);
   M1_2_22_0 : MUX2_X1 port map( A => MR_int_2_22_port, B => MR_int_2_26_port, 
                           S => n35, Z => MR_int_3_22_port);
   M1_2_21_0 : MUX2_X1 port map( A => MR_int_2_21_port, B => MR_int_2_25_port, 
                           S => n35, Z => MR_int_3_21_port);
   M1_2_20_0 : MUX2_X1 port map( A => MR_int_2_20_port, B => MR_int_2_24_port, 
                           S => n35, Z => MR_int_3_20_port);
   M1_2_19_0 : MUX2_X1 port map( A => MR_int_2_19_port, B => MR_int_2_23_port, 
                           S => n35, Z => MR_int_3_19_port);
   M1_2_18_0 : MUX2_X1 port map( A => MR_int_2_18_port, B => MR_int_2_22_port, 
                           S => n35, Z => MR_int_3_18_port);
   M1_2_17_0 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_21_port, 
                           S => n35, Z => MR_int_3_17_port);
   M1_2_16_0 : MUX2_X1 port map( A => MR_int_2_16_port, B => MR_int_2_20_port, 
                           S => n35, Z => MR_int_3_16_port);
   M1_2_15_0 : MUX2_X1 port map( A => MR_int_2_15_port, B => MR_int_2_19_port, 
                           S => n35, Z => MR_int_3_15_port);
   M1_2_14_0 : MUX2_X1 port map( A => MR_int_2_14_port, B => MR_int_2_18_port, 
                           S => n35, Z => MR_int_3_14_port);
   M1_2_13_0 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, 
                           S => n35, Z => MR_int_3_13_port);
   M1_2_12_0 : MUX2_X1 port map( A => MR_int_2_12_port, B => MR_int_2_16_port, 
                           S => n35, Z => MR_int_3_12_port);
   M1_2_11_0 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_15_port, 
                           S => n34, Z => MR_int_3_11_port);
   M1_2_10_0 : MUX2_X1 port map( A => MR_int_2_10_port, B => MR_int_2_14_port, 
                           S => n34, Z => MR_int_3_10_port);
   M1_2_9_0 : MUX2_X1 port map( A => MR_int_2_9_port, B => MR_int_2_13_port, S 
                           => n34, Z => MR_int_3_9_port);
   M1_2_8_0 : MUX2_X1 port map( A => MR_int_2_8_port, B => MR_int_2_12_port, S 
                           => n34, Z => MR_int_3_8_port);
   M1_2_7_0 : MUX2_X1 port map( A => MR_int_2_7_port, B => MR_int_2_11_port, S 
                           => n34, Z => MR_int_3_7_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => n34, Z => MR_int_3_6_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => n34, Z => MR_int_3_5_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => n34, Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           n34, Z => MR_int_3_3_port);
   M1_2_2 : MUX2_X1 port map( A => MR_int_2_2_port, B => MR_int_2_6_port, S => 
                           n34, Z => MR_int_3_2_port);
   M1_2_1 : MUX2_X1 port map( A => MR_int_2_1_port, B => MR_int_2_5_port, S => 
                           n34, Z => MR_int_3_1_port);
   M1_2_0 : MUX2_X1 port map( A => MR_int_2_0_port, B => MR_int_2_4_port, S => 
                           n34, Z => MR_int_3_0_port);
   M1_1_31_0 : MUX2_X1 port map( A => MR_int_1_31_port, B => MR_int_1_1_port, S
                           => n33, Z => MR_int_2_31_port);
   M1_1_30_0 : MUX2_X1 port map( A => MR_int_1_30_port, B => MR_int_1_0_port, S
                           => n33, Z => MR_int_2_30_port);
   M1_1_29_0 : MUX2_X1 port map( A => MR_int_1_29_port, B => MR_int_1_31_port, 
                           S => n33, Z => MR_int_2_29_port);
   M1_1_28_0 : MUX2_X1 port map( A => MR_int_1_28_port, B => MR_int_1_30_port, 
                           S => n33, Z => MR_int_2_28_port);
   M1_1_27_0 : MUX2_X1 port map( A => MR_int_1_27_port, B => MR_int_1_29_port, 
                           S => n33, Z => MR_int_2_27_port);
   M1_1_26_0 : MUX2_X1 port map( A => MR_int_1_26_port, B => MR_int_1_28_port, 
                           S => n33, Z => MR_int_2_26_port);
   M1_1_25_0 : MUX2_X1 port map( A => MR_int_1_25_port, B => MR_int_1_27_port, 
                           S => n33, Z => MR_int_2_25_port);
   M1_1_24_0 : MUX2_X1 port map( A => MR_int_1_24_port, B => MR_int_1_26_port, 
                           S => n33, Z => MR_int_2_24_port);
   M1_1_23_0 : MUX2_X1 port map( A => MR_int_1_23_port, B => MR_int_1_25_port, 
                           S => n32, Z => MR_int_2_23_port);
   M1_1_22_0 : MUX2_X1 port map( A => MR_int_1_22_port, B => MR_int_1_24_port, 
                           S => n32, Z => MR_int_2_22_port);
   M1_1_21_0 : MUX2_X1 port map( A => MR_int_1_21_port, B => MR_int_1_23_port, 
                           S => n32, Z => MR_int_2_21_port);
   M1_1_20_0 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_22_port, 
                           S => n32, Z => MR_int_2_20_port);
   M1_1_19_0 : MUX2_X1 port map( A => MR_int_1_19_port, B => MR_int_1_21_port, 
                           S => n32, Z => MR_int_2_19_port);
   M1_1_18_0 : MUX2_X1 port map( A => MR_int_1_18_port, B => MR_int_1_20_port, 
                           S => n32, Z => MR_int_2_18_port);
   M1_1_17_0 : MUX2_X1 port map( A => MR_int_1_17_port, B => MR_int_1_19_port, 
                           S => n32, Z => MR_int_2_17_port);
   M1_1_16_0 : MUX2_X1 port map( A => MR_int_1_16_port, B => MR_int_1_18_port, 
                           S => n32, Z => MR_int_2_16_port);
   M1_1_15_0 : MUX2_X1 port map( A => MR_int_1_15_port, B => MR_int_1_17_port, 
                           S => n32, Z => MR_int_2_15_port);
   M1_1_14_0 : MUX2_X1 port map( A => MR_int_1_14_port, B => MR_int_1_16_port, 
                           S => n32, Z => MR_int_2_14_port);
   M1_1_13_0 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, 
                           S => n32, Z => MR_int_2_13_port);
   M1_1_12_0 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, 
                           S => n32, Z => MR_int_2_12_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => n31, Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => n31, Z => MR_int_2_10_port);
   M1_1_9_0 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_11_port, S 
                           => n31, Z => MR_int_2_9_port);
   M1_1_8_0 : MUX2_X1 port map( A => MR_int_1_8_port, B => MR_int_1_10_port, S 
                           => n31, Z => MR_int_2_8_port);
   M1_1_7_0 : MUX2_X1 port map( A => MR_int_1_7_port, B => MR_int_1_9_port, S 
                           => n31, Z => MR_int_2_7_port);
   M1_1_6_0 : MUX2_X1 port map( A => MR_int_1_6_port, B => MR_int_1_8_port, S 
                           => n31, Z => MR_int_2_6_port);
   M1_1_5_0 : MUX2_X1 port map( A => MR_int_1_5_port, B => MR_int_1_7_port, S 
                           => n31, Z => MR_int_2_5_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => n31, Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => n31, Z => MR_int_2_3_port);
   M1_1_2_0 : MUX2_X1 port map( A => MR_int_1_2_port, B => MR_int_1_4_port, S 
                           => n31, Z => MR_int_2_2_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => MR_int_1_3_port, S => 
                           n31, Z => MR_int_2_1_port);
   M1_1_0 : MUX2_X1 port map( A => MR_int_1_0_port, B => MR_int_1_2_port, S => 
                           n31, Z => MR_int_2_0_port);
   M1_0_31_0 : MUX2_X1 port map( A => A(31), B => A(0), S => n30, Z => 
                           MR_int_1_31_port);
   M1_0_30_0 : MUX2_X1 port map( A => A(30), B => A(31), S => n30, Z => 
                           MR_int_1_30_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => n30, Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => n30, Z => 
                           MR_int_1_28_port);
   M1_0_27_0 : MUX2_X1 port map( A => A(27), B => A(28), S => n30, Z => 
                           MR_int_1_27_port);
   M1_0_26_0 : MUX2_X1 port map( A => A(26), B => A(27), S => n30, Z => 
                           MR_int_1_26_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => n30, Z => 
                           MR_int_1_25_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => n30, Z => 
                           MR_int_1_24_port);
   M1_0_23_0 : MUX2_X1 port map( A => A(23), B => A(24), S => n29, Z => 
                           MR_int_1_23_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => n29, Z => 
                           MR_int_1_22_port);
   M1_0_21_0 : MUX2_X1 port map( A => A(21), B => A(22), S => n29, Z => 
                           MR_int_1_21_port);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => n29, Z => 
                           MR_int_1_20_port);
   M1_0_19_0 : MUX2_X1 port map( A => A(19), B => A(20), S => n29, Z => 
                           MR_int_1_19_port);
   M1_0_18_0 : MUX2_X1 port map( A => A(18), B => A(19), S => n29, Z => 
                           MR_int_1_18_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => n29, Z => 
                           MR_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => n29, Z => 
                           MR_int_1_16_port);
   M1_0_15_0 : MUX2_X1 port map( A => A(15), B => A(16), S => n29, Z => 
                           MR_int_1_15_port);
   M1_0_14_0 : MUX2_X1 port map( A => A(14), B => A(15), S => n29, Z => 
                           MR_int_1_14_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => n29, Z => 
                           MR_int_1_13_port);
   M1_0_12_0 : MUX2_X1 port map( A => A(12), B => A(13), S => n29, Z => 
                           MR_int_1_12_port);
   M1_0_11_0 : MUX2_X1 port map( A => A(11), B => A(12), S => n28, Z => 
                           MR_int_1_11_port);
   M1_0_10_0 : MUX2_X1 port map( A => A(10), B => A(11), S => n28, Z => 
                           MR_int_1_10_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => n28, Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => n28, Z => 
                           MR_int_1_8_port);
   M1_0_7_0 : MUX2_X1 port map( A => A(7), B => A(8), S => n28, Z => 
                           MR_int_1_7_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => n28, Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => n28, Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => n28, Z => 
                           MR_int_1_4_port);
   M1_0_3_0 : MUX2_X1 port map( A => A(3), B => A(4), S => n28, Z => 
                           MR_int_1_3_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => n28, Z => 
                           MR_int_1_2_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => n28, Z => 
                           MR_int_1_1_port);
   M1_0_0 : MUX2_X1 port map( A => A(0), B => A(1), S => n28, Z => 
                           MR_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(3), Z => n37);
   U3 : BUF_X1 port map( A => SH(3), Z => n38);
   U4 : BUF_X1 port map( A => SH(4), Z => n40);
   U5 : BUF_X1 port map( A => SH(4), Z => n41);
   U6 : BUF_X1 port map( A => SH(3), Z => n39);
   U7 : BUF_X1 port map( A => SH(4), Z => n42);
   U8 : BUF_X1 port map( A => SH(0), Z => n28);
   U9 : BUF_X1 port map( A => SH(0), Z => n29);
   U10 : BUF_X1 port map( A => SH(1), Z => n31);
   U11 : BUF_X1 port map( A => SH(1), Z => n32);
   U12 : BUF_X1 port map( A => SH(2), Z => n34);
   U13 : BUF_X1 port map( A => SH(2), Z => n35);
   U14 : BUF_X1 port map( A => SH(0), Z => n30);
   U15 : BUF_X1 port map( A => SH(1), Z => n33);
   U16 : BUF_X1 port map( A => SH(2), Z => n36);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Shifter_NBIT32_DW_lbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_NBIT32_DW_lbsh_0;

architecture SYN_mx2 of Shifter_NBIT32_DW_lbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n42, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n42, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n42, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n42, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n42, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n42, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n42, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n42, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n41, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n41, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n41, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n41, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n41, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n41, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n41, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n41, Z => B(16));
   M0_4_15 : MUX2_X1 port map( A => ML_int_4_15_port, B => ML_int_4_31_port, S 
                           => n41, Z => B(15));
   M0_4_14 : MUX2_X1 port map( A => ML_int_4_14_port, B => ML_int_4_30_port, S 
                           => n41, Z => B(14));
   M0_4_13 : MUX2_X1 port map( A => ML_int_4_13_port, B => ML_int_4_29_port, S 
                           => n41, Z => B(13));
   M0_4_12 : MUX2_X1 port map( A => ML_int_4_12_port, B => ML_int_4_28_port, S 
                           => n41, Z => B(12));
   M0_4_11 : MUX2_X1 port map( A => ML_int_4_11_port, B => ML_int_4_27_port, S 
                           => n40, Z => B(11));
   M0_4_10 : MUX2_X1 port map( A => ML_int_4_10_port, B => ML_int_4_26_port, S 
                           => n40, Z => B(10));
   M0_4_9 : MUX2_X1 port map( A => ML_int_4_9_port, B => ML_int_4_25_port, S =>
                           n40, Z => B(9));
   M0_4_8 : MUX2_X1 port map( A => ML_int_4_8_port, B => ML_int_4_24_port, S =>
                           n40, Z => B(8));
   M0_4_7 : MUX2_X1 port map( A => ML_int_4_7_port, B => ML_int_4_23_port, S =>
                           n40, Z => B(7));
   M0_4_6 : MUX2_X1 port map( A => ML_int_4_6_port, B => ML_int_4_22_port, S =>
                           n40, Z => B(6));
   M0_4_5 : MUX2_X1 port map( A => ML_int_4_5_port, B => ML_int_4_21_port, S =>
                           n40, Z => B(5));
   M0_4_4 : MUX2_X1 port map( A => ML_int_4_4_port, B => ML_int_4_20_port, S =>
                           n40, Z => B(4));
   M0_4_3 : MUX2_X1 port map( A => ML_int_4_3_port, B => ML_int_4_19_port, S =>
                           n40, Z => B(3));
   M0_4_2 : MUX2_X1 port map( A => ML_int_4_2_port, B => ML_int_4_18_port, S =>
                           n40, Z => B(2));
   M0_4_1 : MUX2_X1 port map( A => ML_int_4_1_port, B => ML_int_4_17_port, S =>
                           n40, Z => B(1));
   M0_4_0 : MUX2_X1 port map( A => ML_int_4_0_port, B => ML_int_4_16_port, S =>
                           n40, Z => B(0));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n39, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n39, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n39, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n39, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n39, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n39, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n39, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n39, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n38, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n38, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n38, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n38, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n38, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n38, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n38, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n38, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n38, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n38, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n38, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n38, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n37, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n37, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n37, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n37, Z => ML_int_4_8_port);
   M0_3_7 : MUX2_X1 port map( A => ML_int_3_7_port, B => ML_int_3_31_port, S =>
                           n37, Z => ML_int_4_7_port);
   M0_3_6 : MUX2_X1 port map( A => ML_int_3_6_port, B => ML_int_3_30_port, S =>
                           n37, Z => ML_int_4_6_port);
   M0_3_5 : MUX2_X1 port map( A => ML_int_3_5_port, B => ML_int_3_29_port, S =>
                           n37, Z => ML_int_4_5_port);
   M0_3_4 : MUX2_X1 port map( A => ML_int_3_4_port, B => ML_int_3_28_port, S =>
                           n37, Z => ML_int_4_4_port);
   M0_3_3 : MUX2_X1 port map( A => ML_int_3_3_port, B => ML_int_3_27_port, S =>
                           n37, Z => ML_int_4_3_port);
   M0_3_2 : MUX2_X1 port map( A => ML_int_3_2_port, B => ML_int_3_26_port, S =>
                           n37, Z => ML_int_4_2_port);
   M0_3_1 : MUX2_X1 port map( A => ML_int_3_1_port, B => ML_int_3_25_port, S =>
                           n37, Z => ML_int_4_1_port);
   M0_3_0 : MUX2_X1 port map( A => ML_int_3_0_port, B => ML_int_3_24_port, S =>
                           n37, Z => ML_int_4_0_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n36, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n36, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n36, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n36, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n36, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n36, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n36, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n36, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n35, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n35, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n35, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n35, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n35, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n35, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n35, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n35, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n35, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n35, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n35, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n35, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n34, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n34, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n34, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n34, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n34, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n34, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n34, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n34, Z => ML_int_3_4_port);
   M0_2_3 : MUX2_X1 port map( A => ML_int_2_3_port, B => ML_int_2_31_port, S =>
                           n34, Z => ML_int_3_3_port);
   M0_2_2 : MUX2_X1 port map( A => ML_int_2_2_port, B => ML_int_2_30_port, S =>
                           n34, Z => ML_int_3_2_port);
   M0_2_1 : MUX2_X1 port map( A => ML_int_2_1_port, B => ML_int_2_29_port, S =>
                           n34, Z => ML_int_3_1_port);
   M0_2_0 : MUX2_X1 port map( A => ML_int_2_0_port, B => ML_int_2_28_port, S =>
                           n34, Z => ML_int_3_0_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n33, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n33, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n33, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n33, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n33, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n33, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n33, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n33, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n32, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n32, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n32, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n32, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n32, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n32, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n32, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n32, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n32, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n32, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n32, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n32, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n31, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n31, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n31, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n31, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n31, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n31, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n31, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n31, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n31, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n31, Z => ML_int_2_2_port);
   M0_1_1 : MUX2_X1 port map( A => ML_int_1_1_port, B => ML_int_1_31_port, S =>
                           n31, Z => ML_int_2_1_port);
   M0_1_0 : MUX2_X1 port map( A => ML_int_1_0_port, B => ML_int_1_30_port, S =>
                           n31, Z => ML_int_2_0_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n30, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n30, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n30, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n30, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n30, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n30, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n30, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n30, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n29, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n29, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n29, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n29, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n29, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n29, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n29, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n29, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n29, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n29, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n29, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n29, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n28, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n28, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n28, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n28, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n28, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n28, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n28, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n28, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n28, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n28, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n28, Z => 
                           ML_int_1_1_port);
   M0_0_0 : MUX2_X1 port map( A => A(0), B => A(31), S => n28, Z => 
                           ML_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(3), Z => n37);
   U3 : BUF_X1 port map( A => SH(3), Z => n38);
   U4 : BUF_X1 port map( A => SH(4), Z => n40);
   U5 : BUF_X1 port map( A => SH(4), Z => n41);
   U6 : BUF_X1 port map( A => SH(3), Z => n39);
   U7 : BUF_X1 port map( A => SH(4), Z => n42);
   U8 : BUF_X1 port map( A => SH(0), Z => n28);
   U9 : BUF_X1 port map( A => SH(0), Z => n29);
   U10 : BUF_X1 port map( A => SH(1), Z => n31);
   U11 : BUF_X1 port map( A => SH(1), Z => n32);
   U12 : BUF_X1 port map( A => SH(2), Z => n34);
   U13 : BUF_X1 port map( A => SH(2), Z => n35);
   U14 : BUF_X1 port map( A => SH(0), Z => n30);
   U15 : BUF_X1 port map( A => SH(1), Z => n33);
   U16 : BUF_X1 port map( A => SH(2), Z => n36);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Shifter_NBIT32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_NBIT32_DW_sra_0;

architecture SYN_mx2 of Shifter_NBIT32_DW_sra_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n73);
   U142 : MUX2_X1 port map( A => A(31), B => A(30), S => n51, Z => n84);
   U3 : NOR2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n51);
   U4 : NOR2_X1 port map( A1 => n183, A2 => SH(1), ZN => n50);
   U5 : NAND2_X1 port map( A1 => n191, A2 => A(31), ZN => n58);
   U6 : INV_X1 port map( A => n38, ZN => n6);
   U7 : INV_X1 port map( A => n191, ZN => n187);
   U8 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n187, A => n5, 
                           ZN => B_9_port);
   U9 : OAI221_X1 port map( B1 => n13, B2 => n3, C1 => n14, C2 => n187, A => 
                           n15, ZN => B_8_port);
   U10 : OAI221_X1 port map( B1 => n115, B2 => n3, C1 => n66, C2 => n187, A => 
                           n116, ZN => B_13_port);
   U11 : OAI221_X1 port map( B1 => n130, B2 => n3, C1 => n67, C2 => n187, A => 
                           n131, ZN => B_12_port);
   U12 : OAI221_X1 port map( B1 => n132, B2 => n3, C1 => n68, C2 => n187, A => 
                           n133, ZN => B_11_port);
   U13 : OAI221_X1 port map( B1 => n148, B2 => n3, C1 => n69, C2 => n187, A => 
                           n149, ZN => B_10_port);
   U14 : NAND2_X1 port map( A1 => n71, A2 => n187, ZN => n38);
   U15 : INV_X1 port map( A => n3, ZN => n41);
   U16 : BUF_X1 port map( A => n186, Z => n190);
   U17 : BUF_X1 port map( A => n185, Z => n188);
   U18 : BUF_X1 port map( A => n185, Z => n189);
   U19 : BUF_X1 port map( A => n186, Z => n191);
   U20 : NOR2_X1 port map( A1 => n184, A2 => SH(3), ZN => n71);
   U21 : INV_X1 port map( A => n54, ZN => n48);
   U22 : INV_X1 port map( A => n56, ZN => n49);
   U23 : INV_X1 port map( A => n50, ZN => n43);
   U24 : INV_X1 port map( A => n51, ZN => n45);
   U25 : NAND2_X1 port map( A1 => n73, A2 => n187, ZN => n3);
   U26 : AOI221_X1 port map( B1 => n84, B2 => n71, C1 => n79, C2 => n73, A => 
                           n74, ZN => n69);
   U27 : AOI221_X1 port map( B1 => n70, B2 => n71, C1 => n72, C2 => n73, A => 
                           n74, ZN => n4);
   U28 : AOI221_X1 port map( B1 => n75, B2 => n71, C1 => n76, C2 => n73, A => 
                           n74, ZN => n14);
   U29 : AOI221_X1 port map( B1 => n77, B2 => n71, C1 => n78, C2 => n73, A => 
                           n74, ZN => n21);
   U30 : AOI221_X1 port map( B1 => n79, B2 => n71, C1 => n80, C2 => n73, A => 
                           n81, ZN => n27);
   U31 : INV_X1 port map( A => n82, ZN => n81);
   U32 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U33 : AOI221_X1 port map( B1 => n72, B2 => n71, C1 => n11, C2 => n73, A => 
                           n86, ZN => n33);
   U34 : INV_X1 port map( A => n87, ZN => n86);
   U35 : AOI21_X1 port map( B1 => n83, B2 => n70, A => n85, ZN => n87);
   U36 : AOI221_X1 port map( B1 => n76, B2 => n71, C1 => n18, C2 => n73, A => 
                           n88, ZN => n36);
   U37 : INV_X1 port map( A => n89, ZN => n88);
   U38 : AOI21_X1 port map( B1 => n83, B2 => n75, A => n85, ZN => n89);
   U39 : AOI221_X1 port map( B1 => n78, B2 => n71, C1 => n25, C2 => n73, A => 
                           n98, ZN => n39);
   U40 : INV_X1 port map( A => n99, ZN => n98);
   U41 : AOI21_X1 port map( B1 => n83, B2 => n77, A => n85, ZN => n99);
   U42 : AOI221_X1 port map( B1 => n80, B2 => n71, C1 => n31, C2 => n73, A => 
                           n102, ZN => n59);
   U43 : INV_X1 port map( A => n103, ZN => n102);
   U44 : AOI22_X1 port map( A1 => n104, A2 => n84, B1 => n83, B2 => n79, ZN => 
                           n103);
   U45 : AOI221_X1 port map( B1 => n11, B2 => n71, C1 => n9, C2 => n73, A => 
                           n105, ZN => n90);
   U46 : INV_X1 port map( A => n106, ZN => n105);
   U47 : AOI22_X1 port map( A1 => n104, A2 => n70, B1 => n83, B2 => n72, ZN => 
                           n106);
   U48 : AOI221_X1 port map( B1 => n18, B2 => n71, C1 => n17, C2 => n73, A => 
                           n162, ZN => n107);
   U49 : INV_X1 port map( A => n163, ZN => n162);
   U50 : AOI22_X1 port map( A1 => n104, A2 => n75, B1 => n83, B2 => n76, ZN => 
                           n163);
   U51 : AOI222_X1 port map( A1 => n6, A2 => n17, B1 => n8, B2 => n18, C1 => 
                           n10, C2 => n76, ZN => n131);
   U52 : AOI222_X1 port map( A1 => n6, A2 => n24, B1 => n8, B2 => n25, C1 => 
                           n10, C2 => n78, ZN => n133);
   U53 : AOI222_X1 port map( A1 => n6, A2 => n30, B1 => n8, B2 => n31, C1 => 
                           n10, C2 => n80, ZN => n149);
   U54 : AOI222_X1 port map( A1 => n6, A2 => n16, B1 => n8, B2 => n17, C1 => 
                           n10, C2 => n18, ZN => n15);
   U55 : AOI222_X1 port map( A1 => n6, A2 => n23, B1 => n8, B2 => n24, C1 => 
                           n10, C2 => n25, ZN => n22);
   U56 : AOI222_X1 port map( A1 => n6, A2 => n29, B1 => n8, B2 => n30, C1 => 
                           n10, C2 => n31, ZN => n28);
   U57 : AOI222_X1 port map( A1 => n6, A2 => n31, B1 => n8, B2 => n80, C1 => 
                           n10, C2 => n79, ZN => n113);
   U58 : AOI222_X1 port map( A1 => n6, A2 => n9, B1 => n8, B2 => n11, C1 => n10
                           , C2 => n72, ZN => n116);
   U59 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10,
                           C2 => n11, ZN => n5);
   U60 : AOI222_X1 port map( A1 => n6, A2 => n12, B1 => n8, B2 => n7, C1 => n10
                           , C2 => n9, ZN => n34);
   U61 : AOI222_X1 port map( A1 => n6, A2 => n19, B1 => n8, B2 => n16, C1 => 
                           n10, C2 => n17, ZN => n37);
   U62 : OAI221_X1 port map( B1 => n20, B2 => n3, C1 => n21, C2 => n187, A => 
                           n22, ZN => B_7_port);
   U63 : OAI221_X1 port map( B1 => n26, B2 => n3, C1 => n27, C2 => n187, A => 
                           n28, ZN => B_6_port);
   U64 : OAI221_X1 port map( B1 => n32, B2 => n3, C1 => n33, C2 => n187, A => 
                           n34, ZN => B_5_port);
   U65 : OAI221_X1 port map( B1 => n35, B2 => n3, C1 => n36, C2 => n187, A => 
                           n37, ZN => B_4_port);
   U66 : OAI221_X1 port map( B1 => n20, B2 => n38, C1 => n39, C2 => n187, A => 
                           n40, ZN => B_3_port);
   U67 : OAI221_X1 port map( B1 => n108, B2 => n38, C1 => n109, C2 => n3, A => 
                           n110, ZN => B_15_port);
   U68 : OAI221_X1 port map( B1 => n112, B2 => n3, C1 => n57, C2 => n187, A => 
                           n113, ZN => B_14_port);
   U69 : OAI221_X1 port map( B1 => n26, B2 => n38, C1 => n59, C2 => n187, A => 
                           n60, ZN => B_2_port);
   U70 : OAI221_X1 port map( B1 => n32, B2 => n38, C1 => n90, C2 => n187, A => 
                           n91, ZN => B_1_port);
   U71 : OAI221_X1 port map( B1 => n35, B2 => n38, C1 => n107, C2 => n187, A =>
                           n156, ZN => B_0_port);
   U72 : OAI21_X1 port map( B1 => n190, B2 => n57, A => n58, ZN => B_30_port);
   U73 : OAI21_X1 port map( B1 => n190, B2 => n66, A => n58, ZN => B_29_port);
   U74 : OAI21_X1 port map( B1 => n190, B2 => n67, A => n58, ZN => B_28_port);
   U75 : OAI21_X1 port map( B1 => n190, B2 => n68, A => n58, ZN => B_27_port);
   U76 : OAI21_X1 port map( B1 => n190, B2 => n69, A => n58, ZN => B_26_port);
   U77 : OAI21_X1 port map( B1 => n189, B2 => n4, A => n58, ZN => B_25_port);
   U78 : OAI21_X1 port map( B1 => n189, B2 => n14, A => n58, ZN => B_24_port);
   U79 : OAI21_X1 port map( B1 => n189, B2 => n21, A => n58, ZN => B_23_port);
   U80 : OAI21_X1 port map( B1 => n189, B2 => n27, A => n58, ZN => B_22_port);
   U81 : OAI21_X1 port map( B1 => n188, B2 => n33, A => n58, ZN => B_21_port);
   U82 : OAI21_X1 port map( B1 => n188, B2 => n36, A => n58, ZN => B_20_port);
   U83 : OAI21_X1 port map( B1 => n188, B2 => n39, A => n58, ZN => B_19_port);
   U84 : OAI21_X1 port map( B1 => n188, B2 => n59, A => n58, ZN => B_18_port);
   U85 : OAI21_X1 port map( B1 => n188, B2 => n90, A => n58, ZN => B_17_port);
   U86 : OAI21_X1 port map( B1 => n189, B2 => n107, A => n58, ZN => B_16_port);
   U87 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n78, A => 
                           n111, ZN => n110);
   U88 : INV_X1 port map( A => n58, ZN => n111);
   U89 : NOR2_X1 port map( A1 => n100, A2 => n184, ZN => n85);
   U90 : AND2_X1 port map( A1 => n159, A2 => n184, ZN => n8);
   U91 : AND2_X1 port map( A1 => SH(3), A2 => n184, ZN => n83);
   U92 : AOI21_X1 port map( B1 => n84, B2 => n73, A => n114, ZN => n57);
   U93 : AOI21_X1 port map( B1 => n70, B2 => n73, A => n114, ZN => n66);
   U94 : AOI21_X1 port map( B1 => n75, B2 => n73, A => n114, ZN => n67);
   U95 : AOI21_X1 port map( B1 => n77, B2 => n73, A => n114, ZN => n68);
   U96 : INV_X1 port map( A => n100, ZN => n74);
   U97 : INV_X1 port map( A => n112, ZN => n30);
   U98 : INV_X1 port map( A => n109, ZN => n24);
   U99 : INV_X1 port map( A => n25, ZN => n108);
   U100 : INV_X1 port map( A => n7, ZN => n115);
   U101 : INV_X1 port map( A => n16, ZN => n130);
   U102 : AND2_X1 port map( A1 => SH(3), A2 => n187, ZN => n159);
   U103 : INV_X1 port map( A => n23, ZN => n132);
   U104 : INV_X1 port map( A => n29, ZN => n148);
   U105 : INV_X1 port map( A => n12, ZN => n2);
   U106 : INV_X1 port map( A => n19, ZN => n13);
   U107 : BUF_X1 port map( A => SH(4), Z => n186);
   U108 : BUF_X1 port map( A => SH(4), Z => n185);
   U109 : OAI221_X1 port map( B1 => n43, B2 => n165, C1 => n45, C2 => n142, A 
                           => n166, ZN => n75);
   U110 : INV_X1 port map( A => A(29), ZN => n165);
   U111 : AOI22_X1 port map( A1 => A(30), A2 => n48, B1 => A(31), B2 => n49, ZN
                           => n166);
   U112 : OAI221_X1 port map( B1 => n43, B2 => n134, C1 => n45, C2 => n135, A 
                           => n136, ZN => n78);
   U113 : AOI22_X1 port map( A1 => A(25), A2 => n48, B1 => A(26), B2 => n49, ZN
                           => n136);
   U114 : OAI221_X1 port map( B1 => n43, B2 => n143, C1 => n45, C2 => n117, A 
                           => n154, ZN => n79);
   U115 : AOI22_X1 port map( A1 => A(28), A2 => n48, B1 => A(29), B2 => n49, ZN
                           => n154);
   U116 : OAI221_X1 port map( B1 => n43, B2 => n117, C1 => n45, C2 => n118, A 
                           => n119, ZN => n72);
   U117 : AOI22_X1 port map( A1 => A(27), A2 => n48, B1 => A(28), B2 => n49, ZN
                           => n119);
   U118 : OAI221_X1 port map( B1 => n43, B2 => n118, C1 => n45, C2 => n134, A 
                           => n164, ZN => n76);
   U119 : AOI22_X1 port map( A1 => A(26), A2 => n48, B1 => A(27), B2 => n49, ZN
                           => n164);
   U120 : OAI221_X1 port map( B1 => n43, B2 => n135, C1 => n45, C2 => n120, A 
                           => n150, ZN => n80);
   U121 : AOI22_X1 port map( A1 => A(24), A2 => n48, B1 => A(25), B2 => n49, ZN
                           => n150);
   U122 : OAI221_X1 port map( B1 => n43, B2 => n120, C1 => n45, C2 => n121, A 
                           => n122, ZN => n11);
   U123 : AOI22_X1 port map( A1 => A(23), A2 => n48, B1 => A(24), B2 => n49, ZN
                           => n122);
   U124 : OAI221_X1 port map( B1 => n43, B2 => n121, C1 => n137, C2 => n45, A 
                           => n168, ZN => n18);
   U125 : AOI22_X1 port map( A1 => A(22), A2 => n48, B1 => A(23), B2 => n49, ZN
                           => n168);
   U126 : OAI221_X1 port map( B1 => n43, B2 => n127, C1 => n45, C2 => n128, A 
                           => n129, ZN => n7);
   U127 : INV_X1 port map( A => A(14), ZN => n127);
   U128 : AOI22_X1 port map( A1 => A(15), A2 => n48, B1 => A(16), B2 => n49, ZN
                           => n129);
   U129 : OAI221_X1 port map( B1 => n43, B2 => n128, C1 => n45, C2 => n145, A 
                           => n161, ZN => n16);
   U130 : AOI22_X1 port map( A1 => A(14), A2 => n48, B1 => A(15), B2 => n49, ZN
                           => n161);
   U131 : OAI221_X1 port map( B1 => n43, B2 => n123, C1 => n45, C2 => n124, A 
                           => n125, ZN => n9);
   U132 : AOI22_X1 port map( A1 => A(19), A2 => n48, B1 => A(20), B2 => n49, ZN
                           => n125);
   U133 : OAI221_X1 port map( B1 => n137, B2 => n43, C1 => n138, C2 => n45, A 
                           => n139, ZN => n25);
   U134 : AOI22_X1 port map( A1 => A(21), A2 => n48, B1 => A(22), B2 => n49, ZN
                           => n139);
   U135 : OAI221_X1 port map( B1 => n138, B2 => n43, C1 => n123, C2 => n45, A 
                           => n151, ZN => n31);
   U136 : AOI22_X1 port map( A1 => A(20), A2 => n48, B1 => A(21), B2 => n49, ZN
                           => n151);
   U137 : OAI221_X1 port map( B1 => n43, B2 => n142, C1 => n45, C2 => n143, A 
                           => n144, ZN => n77);
   U138 : AOI22_X1 port map( A1 => A(29), A2 => n48, B1 => A(30), B2 => n49, ZN
                           => n144);
   U139 : OAI221_X1 port map( B1 => n54, B2 => n123, C1 => n138, C2 => n56, A 
                           => n167, ZN => n17);
   U140 : AOI22_X1 port map( A1 => A(17), A2 => n50, B1 => A(16), B2 => n51, ZN
                           => n167);
   U141 : AOI221_X1 port map( B1 => n50, B2 => A(8), C1 => n51, C2 => A(7), A 
                           => n52, ZN => n20);
   U143 : OAI22_X1 port map( A1 => n53, A2 => n54, B1 => n55, B2 => n56, ZN => 
                           n52);
   U144 : AOI221_X1 port map( B1 => n50, B2 => A(7), C1 => n51, C2 => A(6), A 
                           => n64, ZN => n26);
   U145 : OAI22_X1 port map( A1 => n65, A2 => n54, B1 => n53, B2 => n56, ZN => 
                           n64);
   U146 : AOI221_X1 port map( B1 => n50, B2 => A(6), C1 => n51, C2 => A(5), A 
                           => n96, ZN => n32);
   U147 : OAI22_X1 port map( A1 => n97, A2 => n54, B1 => n65, B2 => n56, ZN => 
                           n96);
   U148 : AOI221_X1 port map( B1 => n50, B2 => A(5), C1 => n51, C2 => A(4), A 
                           => n169, ZN => n35);
   U149 : OAI22_X1 port map( A1 => n170, A2 => n54, B1 => n97, B2 => n56, ZN =>
                           n169);
   U150 : INV_X1 port map( A => A(6), ZN => n170);
   U151 : AOI221_X1 port map( B1 => n50, B2 => A(15), C1 => n51, C2 => A(14), A
                           => n152, ZN => n112);
   U152 : INV_X1 port map( A => n153, ZN => n152);
   U153 : AOI22_X1 port map( A1 => A(16), A2 => n48, B1 => A(17), B2 => n49, ZN
                           => n153);
   U154 : OAI221_X1 port map( B1 => n43, B2 => n145, C1 => n45, C2 => n146, A 
                           => n147, ZN => n23);
   U155 : AOI22_X1 port map( A1 => A(13), A2 => n48, B1 => A(14), B2 => n49, ZN
                           => n147);
   U156 : OAI221_X1 port map( B1 => n43, B2 => n146, C1 => n45, C2 => n55, A =>
                           n155, ZN => n29);
   U157 : AOI22_X1 port map( A1 => A(12), A2 => n48, B1 => A(13), B2 => n49, ZN
                           => n155);
   U158 : OAI221_X1 port map( B1 => n43, B2 => n55, C1 => n45, C2 => n53, A => 
                           n93, ZN => n12);
   U159 : AOI22_X1 port map( A1 => A(11), A2 => n48, B1 => A(12), B2 => n49, ZN
                           => n93);
   U160 : OAI221_X1 port map( B1 => n43, B2 => n53, C1 => n45, C2 => n65, A => 
                           n158, ZN => n19);
   U161 : AOI22_X1 port map( A1 => A(10), A2 => n48, B1 => A(11), B2 => n49, ZN
                           => n158);
   U162 : AOI221_X1 port map( B1 => n50, B2 => A(16), C1 => n51, C2 => A(15), A
                           => n140, ZN => n109);
   U163 : OAI22_X1 port map( A1 => n124, A2 => n54, B1 => n123, B2 => n56, ZN 
                           => n140);
   U164 : AOI222_X1 port map( A1 => n10, A2 => n24, B1 => n41, B2 => n42, C1 =>
                           n8, C2 => n23, ZN => n40);
   U165 : OAI221_X1 port map( B1 => n43, B2 => n44, C1 => n45, C2 => n46, A => 
                           n47, ZN => n42);
   U166 : INV_X1 port map( A => A(4), ZN => n44);
   U167 : AOI22_X1 port map( A1 => A(5), A2 => n48, B1 => A(6), B2 => n49, ZN 
                           => n47);
   U168 : AOI222_X1 port map( A1 => n10, A2 => n30, B1 => n41, B2 => n61, C1 =>
                           n8, C2 => n29, ZN => n60);
   U169 : OAI221_X1 port map( B1 => n43, B2 => n46, C1 => n45, C2 => n62, A => 
                           n63, ZN => n61);
   U170 : AOI22_X1 port map( A1 => A(4), A2 => n48, B1 => A(5), B2 => n49, ZN 
                           => n63);
   U171 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n92, C1 => 
                           n8, C2 => n12, ZN => n91);
   U172 : OAI221_X1 port map( B1 => n43, B2 => n62, C1 => n45, C2 => n94, A => 
                           n95, ZN => n92);
   U173 : INV_X1 port map( A => A(1), ZN => n94);
   U174 : AOI22_X1 port map( A1 => A(3), A2 => n48, B1 => A(4), B2 => n49, ZN 
                           => n95);
   U175 : AOI222_X1 port map( A1 => n10, A2 => n16, B1 => n41, B2 => n157, C1 
                           => n8, C2 => n19, ZN => n156);
   U176 : OAI221_X1 port map( B1 => n54, B2 => n62, C1 => n56, C2 => n46, A => 
                           n160, ZN => n157);
   U177 : AOI22_X1 port map( A1 => A(1), A2 => n50, B1 => A(0), B2 => n51, ZN 
                           => n160);
   U178 : OAI21_X1 port map( B1 => n184, B2 => n141, A => n100, ZN => n114);
   U179 : INV_X1 port map( A => A(31), ZN => n141);
   U180 : NAND2_X1 port map( A1 => SH(1), A2 => n183, ZN => n54);
   U181 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n56);
   U182 : AND2_X1 port map( A1 => SH(2), A2 => n159, ZN => n10);
   U183 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n100);
   U184 : INV_X1 port map( A => n126, ZN => n70);
   U185 : AOI222_X1 port map( A1 => n51, A2 => A(29), B1 => n50, B2 => A(30), 
                           C1 => SH(1), C2 => A(31), ZN => n126);
   U186 : INV_X1 port map( A => A(9), ZN => n53);
   U187 : INV_X1 port map( A => A(18), ZN => n123);
   U188 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n104);
   U189 : INV_X1 port map( A => A(3), ZN => n46);
   U190 : INV_X1 port map( A => A(8), ZN => n65);
   U191 : INV_X1 port map( A => A(10), ZN => n55);
   U192 : INV_X1 port map( A => A(2), ZN => n62);
   U193 : INV_X1 port map( A => A(19), ZN => n138);
   U194 : INV_X1 port map( A => A(20), ZN => n137);
   U195 : INV_X1 port map( A => A(17), ZN => n124);
   U196 : INV_X1 port map( A => A(11), ZN => n146);
   U197 : INV_X1 port map( A => A(12), ZN => n145);
   U198 : INV_X1 port map( A => A(13), ZN => n128);
   U199 : INV_X1 port map( A => A(28), ZN => n142);
   U200 : INV_X1 port map( A => A(27), ZN => n143);
   U201 : INV_X1 port map( A => A(26), ZN => n117);
   U202 : INV_X1 port map( A => A(25), ZN => n118);
   U203 : INV_X1 port map( A => A(24), ZN => n134);
   U204 : INV_X1 port map( A => A(23), ZN => n135);
   U205 : INV_X1 port map( A => A(22), ZN => n120);
   U206 : INV_X1 port map( A => A(21), ZN => n121);
   U207 : INV_X1 port map( A => A(7), ZN => n97);
   U208 : INV_X1 port map( A => SH(0), ZN => n183);
   U209 : INV_X1 port map( A => SH(2), ZN => n184);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Shifter_NBIT32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end Shifter_NBIT32_DW_rash_0;

architecture SYN_mx2 of Shifter_NBIT32_DW_rash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n149, n150, n151, 
      n152, n154, n155, n156, n157, n158, n159, n160, n161, n163, n164, n165, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191 : 
      std_logic;

begin
   
   U102 : MUX2_X1 port map( A => n75, B => n58, S => SH(2), Z => n89);
   U3 : NOR2_X1 port map( A1 => n182, A2 => n183, ZN => n73);
   U4 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n44);
   U5 : INV_X1 port map( A => n3, ZN => n41);
   U6 : NAND2_X1 port map( A1 => n72, A2 => n191, ZN => n3);
   U7 : INV_X1 port map( A => n188, ZN => n191);
   U8 : INV_X1 port map( A => n38, ZN => n6);
   U9 : INV_X1 port map( A => n164, ZN => n52);
   U10 : NAND2_X1 port map( A1 => n73, A2 => n191, ZN => n38);
   U11 : NOR2_X1 port map( A1 => n191, A2 => n124, ZN => n99);
   U12 : INV_X1 port map( A => n124, ZN => n72);
   U13 : NOR2_X1 port map( A1 => n184, A2 => n185, ZN => n147);
   U14 : BUF_X1 port map( A => n190, Z => n185);
   U15 : BUF_X1 port map( A => n190, Z => n186);
   U16 : BUF_X1 port map( A => n189, Z => n187);
   U17 : BUF_X1 port map( A => n189, Z => n188);
   U18 : OAI222_X1 port map( A1 => n55, A2 => n109, B1 => n163, B2 => n110, C1 
                           => n57, C2 => n111, ZN => n67);
   U19 : INV_X1 port map( A => n50, ZN => n57);
   U20 : OAI22_X1 port map( A1 => n57, A2 => n109, B1 => n55, B2 => n110, ZN =>
                           n59);
   U21 : AOI222_X1 port map( A1 => n23, A2 => n72, B1 => n77, B2 => n73, C1 => 
                           n89, C2 => n183, ZN => n39);
   U22 : AOI222_X1 port map( A1 => n75, A2 => n73, B1 => n58, B2 => n76, C1 => 
                           n77, C2 => n72, ZN => n19);
   U23 : AOI222_X1 port map( A1 => n78, A2 => n73, B1 => n59, B2 => n76, C1 => 
                           n79, C2 => n72, ZN => n25);
   U24 : AOI222_X1 port map( A1 => n71, A2 => n73, B1 => n67, B2 => n76, C1 => 
                           n11, C2 => n72, ZN => n31);
   U25 : AOI222_X1 port map( A1 => n74, A2 => n73, B1 => n68, B2 => n76, C1 => 
                           n17, C2 => n72, ZN => n35);
   U26 : INV_X1 port map( A => n49, ZN => n55);
   U27 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n29, C2 => n72, A => 
                           n90, ZN => n60);
   U28 : INV_X1 port map( A => n91, ZN => n90);
   U29 : AOI22_X1 port map( A1 => n92, A2 => n59, B1 => n76, B2 => n78, ZN => 
                           n91);
   U30 : AOI221_X1 port map( B1 => n11, B2 => n73, C1 => n9, C2 => n72, A => 
                           n93, ZN => n80);
   U31 : INV_X1 port map( A => n94, ZN => n93);
   U32 : AOI22_X1 port map( A1 => n92, A2 => n67, B1 => n76, B2 => n71, ZN => 
                           n94);
   U33 : AOI221_X1 port map( B1 => n17, B2 => n73, C1 => n16, C2 => n72, A => 
                           n154, ZN => n95);
   U34 : INV_X1 port map( A => n155, ZN => n154);
   U35 : AOI22_X1 port map( A1 => n92, A2 => n68, B1 => n76, B2 => n74, ZN => 
                           n155);
   U36 : AOI222_X1 port map( A1 => n10, A2 => n71, B1 => n99, B2 => n67, C1 => 
                           n8, C2 => n11, ZN => n105);
   U37 : AOI222_X1 port map( A1 => n6, A2 => n28, B1 => n8, B2 => n29, C1 => 
                           n10, C2 => n79, ZN => n138);
   U38 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10,
                           C2 => n11, ZN => n5);
   U39 : AOI222_X1 port map( A1 => n6, A2 => n15, B1 => n8, B2 => n16, C1 => 
                           n10, C2 => n17, ZN => n14);
   U40 : AOI222_X1 port map( A1 => n6, A2 => n27, B1 => n8, B2 => n28, C1 => 
                           n10, C2 => n29, ZN => n26);
   U41 : AOI222_X1 port map( A1 => n6, A2 => n33, B1 => n8, B2 => n7, C1 => n10
                           , C2 => n9, ZN => n32);
   U42 : AOI222_X1 port map( A1 => n6, A2 => n37, B1 => n8, B2 => n15, C1 => 
                           n10, C2 => n16, ZN => n36);
   U43 : AOI222_X1 port map( A1 => n10, A2 => n78, B1 => n99, B2 => n59, C1 => 
                           n8, C2 => n79, ZN => n102);
   U44 : AOI222_X1 port map( A1 => n6, A2 => n21, B1 => n8, B2 => n22, C1 => 
                           n10, C2 => n23, ZN => n20);
   U45 : AOI222_X1 port map( A1 => n10, A2 => n75, B1 => n99, B2 => n58, C1 => 
                           n8, C2 => n77, ZN => n98);
   U46 : INV_X1 port map( A => n44, ZN => n51);
   U47 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n191, A => n5,
                           ZN => B(9));
   U48 : OAI221_X1 port map( B1 => n12, B2 => n3, C1 => n13, C2 => n191, A => 
                           n14, ZN => B(8));
   U49 : OAI221_X1 port map( B1 => n18, B2 => n3, C1 => n19, C2 => n191, A => 
                           n20, ZN => B(7));
   U50 : OAI221_X1 port map( B1 => n24, B2 => n3, C1 => n25, C2 => n191, A => 
                           n26, ZN => B(6));
   U51 : OAI221_X1 port map( B1 => n30, B2 => n3, C1 => n31, C2 => n191, A => 
                           n32, ZN => B(5));
   U52 : OAI221_X1 port map( B1 => n34, B2 => n3, C1 => n35, C2 => n191, A => 
                           n36, ZN => B(4));
   U53 : OAI221_X1 port map( B1 => n18, B2 => n38, C1 => n39, C2 => n191, A => 
                           n40, ZN => B(3));
   U54 : AND2_X1 port map( A1 => n41, A2 => n58, ZN => B(31));
   U55 : OAI221_X1 port map( B1 => n96, B2 => n38, C1 => n97, C2 => n3, A => 
                           n98, ZN => B(15));
   U56 : OAI221_X1 port map( B1 => n100, B2 => n38, C1 => n101, C2 => n3, A => 
                           n102, ZN => B(14));
   U57 : OAI221_X1 port map( B1 => n103, B2 => n38, C1 => n104, C2 => n3, A => 
                           n105, ZN => B(13));
   U58 : INV_X1 port map( A => n121, ZN => B(12));
   U59 : OAI221_X1 port map( B1 => n97, B2 => n38, C1 => n43, C2 => n3, A => 
                           n125, ZN => B(11));
   U60 : OAI221_X1 port map( B1 => n63, B2 => n3, C1 => n70, C2 => n191, A => 
                           n138, ZN => B(10));
   U61 : OAI221_X1 port map( B1 => n24, B2 => n38, C1 => n60, C2 => n191, A => 
                           n61, ZN => B(2));
   U62 : OAI221_X1 port map( B1 => n30, B2 => n38, C1 => n80, C2 => n191, A => 
                           n81, ZN => B(1));
   U63 : AND2_X1 port map( A1 => n59, A2 => n41, ZN => B(30));
   U64 : AND2_X1 port map( A1 => n67, A2 => n41, ZN => B(29));
   U65 : AND2_X1 port map( A1 => n68, A2 => n41, ZN => B(28));
   U66 : NOR3_X1 port map( A1 => n69, A2 => n185, A3 => n183, ZN => B(27));
   U67 : NOR2_X1 port map( A1 => n187, A2 => n70, ZN => B(26));
   U68 : NOR2_X1 port map( A1 => n187, A2 => n4, ZN => B(25));
   U69 : NOR2_X1 port map( A1 => n186, A2 => n13, ZN => B(24));
   U70 : NOR2_X1 port map( A1 => n187, A2 => n19, ZN => B(23));
   U71 : NOR2_X1 port map( A1 => n185, A2 => n25, ZN => B(22));
   U72 : NOR2_X1 port map( A1 => n186, A2 => n31, ZN => B(21));
   U73 : NOR2_X1 port map( A1 => n186, A2 => n35, ZN => B(20));
   U74 : NOR2_X1 port map( A1 => n185, A2 => n39, ZN => B(19));
   U75 : NOR2_X1 port map( A1 => n186, A2 => n60, ZN => B(18));
   U76 : NOR2_X1 port map( A1 => n188, A2 => n80, ZN => B(17));
   U77 : NOR2_X1 port map( A1 => n187, A2 => n95, ZN => B(16));
   U78 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n23, A => 
                           n126, ZN => n125);
   U79 : NOR3_X1 port map( A1 => n191, A2 => n183, A3 => n69, ZN => n126);
   U80 : AOI221_X1 port map( B1 => n16, B2 => n6, C1 => n15, C2 => n41, A => 
                           n122, ZN => n121);
   U81 : INV_X1 port map( A => n123, ZN => n122);
   U82 : AOI222_X1 port map( A1 => n10, A2 => n74, B1 => n99, B2 => n68, C1 => 
                           n8, C2 => n17, ZN => n123);
   U83 : AND2_X1 port map( A1 => n147, A2 => n182, ZN => n8);
   U84 : NOR2_X1 port map( A1 => n110, A2 => n57, ZN => n58);
   U85 : AOI22_X1 port map( A1 => n78, A2 => n72, B1 => n59, B2 => n73, ZN => 
                           n70);
   U86 : AOI22_X1 port map( A1 => n71, A2 => n72, B1 => n67, B2 => n73, ZN => 
                           n4);
   U87 : AOI22_X1 port map( A1 => n74, A2 => n72, B1 => n68, B2 => n73, ZN => 
                           n13);
   U88 : NOR2_X1 port map( A1 => n182, A2 => n184, ZN => n92);
   U89 : BUF_X1 port map( A => n46, Z => n163);
   U90 : BUF_X1 port map( A => n46, Z => n164);
   U91 : BUF_X1 port map( A => n46, Z => n165);
   U92 : INV_X1 port map( A => SH(3), ZN => n184);
   U93 : NAND2_X1 port map( A1 => n182, A2 => n184, ZN => n124);
   U94 : INV_X1 port map( A => n63, ZN => n27);
   U95 : INV_X1 port map( A => n2, ZN => n33);
   U96 : INV_X1 port map( A => n12, ZN => n37);
   U97 : INV_X1 port map( A => n22, ZN => n97);
   U98 : INV_X1 port map( A => n43, ZN => n21);
   U99 : INV_X1 port map( A => n23, ZN => n96);
   U100 : INV_X1 port map( A => n29, ZN => n100);
   U101 : INV_X1 port map( A => n9, ZN => n103);
   U103 : INV_X1 port map( A => n28, ZN => n101);
   U104 : INV_X1 port map( A => n7, ZN => n104);
   U105 : INV_X1 port map( A => n89, ZN => n69);
   U106 : BUF_X1 port map( A => SH(4), Z => n190);
   U107 : BUF_X1 port map( A => SH(4), Z => n189);
   U108 : NOR2_X2 port map( A1 => n181, A2 => SH(1), ZN => n49);
   U109 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n50);
   U110 : OAI221_X1 port map( B1 => n44, B2 => n110, C1 => n164, C2 => n109, A 
                           => n157, ZN => n68);
   U111 : AOI22_X1 port map( A1 => A(29), A2 => n49, B1 => A(28), B2 => n50, ZN
                           => n157);
   U112 : NOR2_X1 port map( A1 => n184, A2 => SH(2), ZN => n76);
   U113 : OAI221_X1 port map( B1 => n118, B2 => n55, C1 => n119, C2 => n57, A 
                           => n128, ZN => n23);
   U114 : AOI22_X1 port map( A1 => A(22), A2 => n51, B1 => A(21), B2 => n52, ZN
                           => n128);
   U115 : OAI221_X1 port map( B1 => n119, B2 => n55, C1 => n135, C2 => n57, A 
                           => n140, ZN => n29);
   U116 : AOI22_X1 port map( A1 => A(21), A2 => n51, B1 => n52, B2 => A(20), ZN
                           => n140);
   U117 : OAI221_X1 port map( B1 => n44, B2 => n118, C1 => n164, C2 => n119, A 
                           => n120, ZN => n9);
   U118 : AOI22_X1 port map( A1 => A(18), A2 => n49, B1 => A(17), B2 => n50, ZN
                           => n120);
   U119 : OAI221_X1 port map( B1 => n44, B2 => n119, C1 => n164, C2 => n135, A 
                           => n158, ZN => n16);
   U120 : AOI22_X1 port map( A1 => A(17), A2 => n49, B1 => A(16), B2 => n50, ZN
                           => n158);
   U121 : OAI221_X1 port map( B1 => n44, B2 => n136, C1 => n165, C2 => n115, A 
                           => n141, ZN => n28);
   U122 : AOI22_X1 port map( A1 => A(15), A2 => n49, B1 => A(14), B2 => n50, ZN
                           => n141);
   U123 : OAI221_X1 port map( B1 => n44, B2 => n115, C1 => n163, C2 => n116, A 
                           => n117, ZN => n7);
   U124 : AOI22_X1 port map( A1 => A(14), A2 => n49, B1 => A(13), B2 => n50, ZN
                           => n117);
   U125 : OAI221_X1 port map( B1 => n44, B2 => n116, C1 => n163, C2 => n151, A 
                           => n152, ZN => n15);
   U126 : INV_X1 port map( A => A(14), ZN => n151);
   U127 : AOI22_X1 port map( A1 => A(13), A2 => n49, B1 => A(12), B2 => n50, ZN
                           => n152);
   U128 : OAI221_X1 port map( B1 => n44, B2 => n111, C1 => n163, C2 => n112, A 
                           => n142, ZN => n78);
   U129 : AOI22_X1 port map( A1 => A(27), A2 => n49, B1 => A(26), B2 => n50, ZN
                           => n142);
   U130 : OAI221_X1 port map( B1 => n44, B2 => n112, C1 => n163, C2 => n113, A 
                           => n114, ZN => n71);
   U131 : AOI22_X1 port map( A1 => A(26), A2 => n49, B1 => A(25), B2 => n50, ZN
                           => n114);
   U132 : OAI221_X1 port map( B1 => n44, B2 => n113, C1 => n164, C2 => n129, A 
                           => n156, ZN => n74);
   U133 : AOI22_X1 port map( A1 => A(25), A2 => n49, B1 => A(24), B2 => n50, ZN
                           => n156);
   U134 : OAI221_X1 port map( B1 => n55, B2 => n159, C1 => n118, C2 => n57, A 
                           => n160, ZN => n17);
   U135 : INV_X1 port map( A => A(21), ZN => n159);
   U136 : AOI22_X1 port map( A1 => A(23), A2 => n51, B1 => A(22), B2 => n52, ZN
                           => n160);
   U137 : OAI221_X1 port map( B1 => n44, B2 => n130, C1 => n165, C2 => n106, A 
                           => n139, ZN => n79);
   U138 : AOI22_X1 port map( A1 => A(23), A2 => n49, B1 => A(22), B2 => n50, ZN
                           => n139);
   U139 : OAI221_X1 port map( B1 => n44, B2 => n106, C1 => n163, C2 => n107, A 
                           => n108, ZN => n11);
   U140 : INV_X1 port map( A => A(23), ZN => n107);
   U141 : AOI22_X1 port map( A1 => A(22), A2 => n49, B1 => A(21), B2 => n50, ZN
                           => n108);
   U142 : OAI221_X1 port map( B1 => n44, B2 => n129, C1 => n164, C2 => n130, A 
                           => n131, ZN => n77);
   U143 : AOI22_X1 port map( A1 => A(24), A2 => n49, B1 => A(23), B2 => n50, ZN
                           => n131);
   U144 : AOI221_X1 port map( B1 => n51, B2 => A(10), C1 => n52, C2 => A(9), A 
                           => n53, ZN => n18);
   U145 : OAI22_X1 port map( A1 => n54, A2 => n55, B1 => n56, B2 => n57, ZN => 
                           n53);
   U146 : AOI221_X1 port map( B1 => n51, B2 => A(9), C1 => n52, C2 => A(8), A 
                           => n66, ZN => n24);
   U147 : OAI22_X1 port map( A1 => n56, A2 => n55, B1 => n45, B2 => n57, ZN => 
                           n66);
   U148 : AOI221_X1 port map( B1 => n51, B2 => A(8), C1 => n52, C2 => A(7), A 
                           => n88, ZN => n30);
   U149 : OAI22_X1 port map( A1 => n45, A2 => n55, B1 => n47, B2 => n57, ZN => 
                           n88);
   U150 : AOI221_X1 port map( B1 => n51, B2 => A(7), C1 => n52, C2 => A(6), A 
                           => n161, ZN => n34);
   U151 : OAI22_X1 port map( A1 => n47, A2 => n55, B1 => n64, B2 => n57, ZN => 
                           n161);
   U152 : AOI221_X1 port map( B1 => n51, B2 => A(13), C1 => n52, C2 => A(12), A
                           => n143, ZN => n63);
   U153 : OAI22_X1 port map( A1 => n134, A2 => n55, B1 => n84, B2 => n57, ZN =>
                           n143);
   U154 : AOI221_X1 port map( B1 => n51, B2 => A(12), C1 => n52, C2 => A(11), A
                           => n83, ZN => n2);
   U155 : OAI22_X1 port map( A1 => n84, A2 => n55, B1 => n85, B2 => n57, ZN => 
                           n83);
   U156 : AOI221_X1 port map( B1 => n51, B2 => A(11), C1 => n52, C2 => A(10), A
                           => n146, ZN => n12);
   U157 : OAI22_X1 port map( A1 => n85, A2 => n55, B1 => n54, B2 => n57, ZN => 
                           n146);
   U158 : OAI221_X1 port map( B1 => n44, B2 => n135, C1 => n165, C2 => n136, A 
                           => n137, ZN => n22);
   U159 : AOI22_X1 port map( A1 => A(16), A2 => n49, B1 => A(15), B2 => n50, ZN
                           => n137);
   U160 : AOI221_X1 port map( B1 => n51, B2 => A(14), C1 => n52, C2 => A(13), A
                           => n132, ZN => n43);
   U161 : OAI22_X1 port map( A1 => n133, A2 => n55, B1 => n134, B2 => n57, ZN 
                           => n132);
   U162 : INV_X1 port map( A => A(12), ZN => n133);
   U163 : AOI222_X1 port map( A1 => n10, A2 => n22, B1 => n41, B2 => n42, C1 =>
                           n8, C2 => n21, ZN => n40);
   U164 : OAI221_X1 port map( B1 => n44, B2 => n45, C1 => n165, C2 => n47, A =>
                           n48, ZN => n42);
   U165 : AOI22_X1 port map( A1 => A(4), A2 => n49, B1 => A(3), B2 => n50, ZN 
                           => n48);
   U166 : AOI222_X1 port map( A1 => n10, A2 => n28, B1 => n41, B2 => n62, C1 =>
                           n8, C2 => n27, ZN => n61);
   U167 : OAI221_X1 port map( B1 => n44, B2 => n47, C1 => n165, C2 => n64, A =>
                           n65, ZN => n62);
   U168 : AOI22_X1 port map( A1 => A(3), A2 => n49, B1 => A(2), B2 => n50, ZN 
                           => n65);
   U169 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n82, C1 => 
                           n8, C2 => n33, ZN => n81);
   U170 : OAI221_X1 port map( B1 => n44, B2 => n64, C1 => n165, C2 => n86, A =>
                           n87, ZN => n82);
   U171 : AOI22_X1 port map( A1 => A(2), A2 => n49, B1 => A(1), B2 => n50, ZN 
                           => n87);
   U172 : OAI221_X1 port map( B1 => n34, B2 => n38, C1 => n95, C2 => n191, A =>
                           n144, ZN => B(0));
   U173 : AOI222_X1 port map( A1 => n10, A2 => n15, B1 => n41, B2 => n145, C1 
                           => n8, C2 => n37, ZN => n144);
   U174 : OAI221_X1 port map( B1 => n44, B2 => n109, C1 => n164, C2 => n111, A 
                           => n127, ZN => n75);
   U175 : AOI22_X1 port map( A1 => A(28), A2 => n49, B1 => A(27), B2 => n50, ZN
                           => n127);
   U176 : OAI221_X1 port map( B1 => n44, B2 => n86, C1 => n163, C2 => n149, A 
                           => n150, ZN => n145);
   U177 : INV_X1 port map( A => A(2), ZN => n149);
   U178 : AOI22_X1 port map( A1 => A(1), A2 => n49, B1 => A(0), B2 => n50, ZN 
                           => n150);
   U179 : AND2_X1 port map( A1 => SH(2), A2 => n147, ZN => n10);
   U180 : INV_X1 port map( A => A(19), ZN => n119);
   U181 : INV_X1 port map( A => A(30), ZN => n109);
   U182 : INV_X1 port map( A => A(31), ZN => n110);
   U183 : INV_X1 port map( A => A(5), ZN => n47);
   U184 : INV_X1 port map( A => A(20), ZN => n118);
   U185 : INV_X1 port map( A => A(4), ZN => n64);
   U186 : INV_X1 port map( A => A(29), ZN => n111);
   U187 : INV_X1 port map( A => A(6), ZN => n45);
   U188 : INV_X1 port map( A => A(18), ZN => n135);
   U189 : NAND2_X1 port map( A1 => SH(1), A2 => n181, ZN => n46);
   U190 : INV_X1 port map( A => A(17), ZN => n136);
   U191 : INV_X1 port map( A => A(16), ZN => n115);
   U192 : INV_X1 port map( A => A(15), ZN => n116);
   U193 : INV_X1 port map( A => A(3), ZN => n86);
   U194 : INV_X1 port map( A => A(28), ZN => n112);
   U195 : INV_X1 port map( A => A(27), ZN => n113);
   U196 : INV_X1 port map( A => A(26), ZN => n129);
   U197 : INV_X1 port map( A => A(25), ZN => n130);
   U198 : INV_X1 port map( A => A(24), ZN => n106);
   U199 : INV_X1 port map( A => A(11), ZN => n134);
   U200 : INV_X1 port map( A => A(10), ZN => n84);
   U201 : INV_X1 port map( A => A(9), ZN => n85);
   U202 : INV_X1 port map( A => A(8), ZN => n54);
   U203 : INV_X1 port map( A => A(7), ZN => n56);
   U204 : INV_X1 port map( A => SH(0), ZN => n181);
   U205 : INV_X1 port map( A => SH(2), ZN => n182);
   U206 : INV_X1 port map( A => n184, ZN => n183);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Shifter_NBIT32_DW_sla_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_NBIT32_DW_sla_0;

architecture SYN_mx2 of Shifter_NBIT32_DW_sla_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78
      , n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n170, n171, n172, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   B <= ( B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, A(0) );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n75);
   U142 : MUX2_X1 port map( A => A(1), B => A(0), S => n34, Z => n79);
   U3 : NAND2_X1 port map( A1 => n195, A2 => A(0), ZN => n3);
   U4 : NAND2_X1 port map( A1 => SH(0), A2 => n187, ZN => n33);
   U5 : INV_X1 port map( A => n11, ZN => n58);
   U6 : INV_X1 port map( A => n195, ZN => n191);
   U7 : INV_X1 port map( A => n34, ZN => n26);
   U8 : NAND2_X1 port map( A1 => n73, A2 => n191, ZN => n11);
   U9 : INV_X1 port map( A => n55, ZN => n16);
   U10 : BUF_X1 port map( A => n190, Z => n194);
   U11 : BUF_X1 port map( A => n189, Z => n192);
   U12 : BUF_X1 port map( A => n189, Z => n193);
   U13 : BUF_X1 port map( A => n190, Z => n195);
   U14 : NOR2_X1 port map( A1 => n188, A2 => SH(3), ZN => n73);
   U15 : INV_X1 port map( A => n20, ZN => n37);
   U16 : INV_X1 port map( A => n22, ZN => n38);
   U17 : OAI222_X1 port map( A1 => n34, A2 => n153, B1 => n154, B2 => n33, C1 
                           => n124, C2 => n187, ZN => n101);
   U18 : NAND2_X1 port map( A1 => n75, A2 => n191, ZN => n55);
   U19 : INV_X1 port map( A => n33, ZN => n25);
   U20 : AOI221_X1 port map( B1 => n86, B2 => n73, C1 => n87, C2 => n75, A => 
                           n88, ZN => n4);
   U21 : AOI221_X1 port map( B1 => n94, B2 => n73, C1 => n95, C2 => n75, A => 
                           n88, ZN => n5);
   U22 : AOI221_X1 port map( B1 => n101, B2 => n73, C1 => n102, C2 => n75, A =>
                           n88, ZN => n6);
   U23 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n72, C2 => n75, A => 
                           n88, ZN => n7);
   U24 : AOI221_X1 port map( B1 => n92, B2 => n73, C1 => n59, C2 => n75, A => 
                           n134, ZN => n12);
   U25 : INV_X1 port map( A => n135, ZN => n134);
   U26 : AOI22_X1 port map( A1 => n136, A2 => n94, B1 => n78, B2 => n95, ZN => 
                           n135);
   U27 : AOI221_X1 port map( B1 => n99, B2 => n73, C1 => n65, C2 => n75, A => 
                           n138, ZN => n28);
   U28 : INV_X1 port map( A => n139, ZN => n138);
   U29 : AOI22_X1 port map( A1 => n136, A2 => n101, B1 => n78, B2 => n102, ZN 
                           => n139);
   U30 : AOI221_X1 port map( B1 => n74, B2 => n73, C1 => n70, C2 => n75, A => 
                           n141, ZN => n41);
   U31 : INV_X1 port map( A => n142, ZN => n141);
   U32 : AOI22_X1 port map( A1 => n136, A2 => n79, B1 => n78, B2 => n72, ZN => 
                           n142);
   U33 : AOI221_X1 port map( B1 => n87, B2 => n73, C1 => n84, C2 => n75, A => 
                           n151, ZN => n48);
   U34 : INV_X1 port map( A => n152, ZN => n151);
   U35 : AOI21_X1 port map( B1 => n78, B2 => n86, A => n80, ZN => n152);
   U36 : AOI221_X1 port map( B1 => n95, B2 => n73, C1 => n92, C2 => n75, A => 
                           n160, ZN => n56);
   U37 : INV_X1 port map( A => n161, ZN => n160);
   U38 : AOI21_X1 port map( B1 => n78, B2 => n94, A => n80, ZN => n161);
   U39 : AOI221_X1 port map( B1 => n102, B2 => n73, C1 => n99, C2 => n75, A => 
                           n167, ZN => n63);
   U40 : INV_X1 port map( A => n168, ZN => n167);
   U41 : AOI21_X1 port map( B1 => n78, B2 => n101, A => n80, ZN => n168);
   U42 : AOI221_X1 port map( B1 => n72, B2 => n73, C1 => n74, C2 => n75, A => 
                           n76, ZN => n2);
   U43 : INV_X1 port map( A => n77, ZN => n76);
   U44 : AOI21_X1 port map( B1 => n78, B2 => n79, A => n80, ZN => n77);
   U45 : AOI222_X1 port map( A1 => n58, A2 => n15, B1 => n18, B2 => n59, C1 => 
                           n14, C2 => n92, ZN => n91);
   U46 : AOI222_X1 port map( A1 => n58, A2 => n30, B1 => n18, B2 => n65, C1 => 
                           n14, C2 => n99, ZN => n98);
   U47 : AOI222_X1 port map( A1 => n58, A2 => n43, B1 => n18, B2 => n70, C1 => 
                           n14, C2 => n74, ZN => n105);
   U48 : AOI222_X1 port map( A1 => n58, A2 => n50, B1 => n18, B2 => n84, C1 => 
                           n14, C2 => n87, ZN => n111);
   U49 : AOI222_X1 port map( A1 => n58, A2 => n59, B1 => n18, B2 => n92, C1 => 
                           n14, C2 => n95, ZN => n117);
   U50 : AOI222_X1 port map( A1 => n58, A2 => n65, B1 => n18, B2 => n99, C1 => 
                           n14, C2 => n102, ZN => n120);
   U51 : AOI222_X1 port map( A1 => n58, A2 => n70, B1 => n18, B2 => n74, C1 => 
                           n14, C2 => n72, ZN => n123);
   U52 : AOI222_X1 port map( A1 => n58, A2 => n19, B1 => n18, B2 => n15, C1 => 
                           n14, C2 => n59, ZN => n57);
   U53 : AOI222_X1 port map( A1 => n58, A2 => n32, B1 => n18, B2 => n30, C1 => 
                           n14, C2 => n65, ZN => n64);
   U54 : AOI222_X1 port map( A1 => n58, A2 => n45, B1 => n18, B2 => n43, C1 => 
                           n14, C2 => n70, ZN => n69);
   U55 : AOI222_X1 port map( A1 => n58, A2 => n52, B1 => n18, B2 => n50, C1 => 
                           n14, C2 => n84, ZN => n83);
   U56 : OAI21_X1 port map( B1 => n194, B2 => n2, A => n3, ZN => B_9_port);
   U57 : OAI21_X1 port map( B1 => n194, B2 => n4, A => n3, ZN => B_8_port);
   U58 : OAI21_X1 port map( B1 => n194, B2 => n5, A => n3, ZN => B_7_port);
   U59 : OAI21_X1 port map( B1 => n194, B2 => n6, A => n3, ZN => B_6_port);
   U60 : OAI21_X1 port map( B1 => n194, B2 => n7, A => n3, ZN => B_5_port);
   U61 : OAI21_X1 port map( B1 => n192, B2 => n8, A => n3, ZN => B_4_port);
   U62 : OAI21_X1 port map( B1 => n192, B2 => n9, A => n3, ZN => B_3_port);
   U63 : OAI221_X1 port map( B1 => n10, B2 => n11, C1 => n12, C2 => n191, A => 
                           n13, ZN => B_31_port);
   U64 : OAI21_X1 port map( B1 => n193, B2 => n12, A => n3, ZN => B_15_port);
   U65 : OAI21_X1 port map( B1 => n193, B2 => n28, A => n3, ZN => B_14_port);
   U66 : OAI21_X1 port map( B1 => n192, B2 => n41, A => n3, ZN => B_13_port);
   U67 : OAI21_X1 port map( B1 => n193, B2 => n48, A => n3, ZN => B_12_port);
   U68 : OAI21_X1 port map( B1 => n193, B2 => n56, A => n3, ZN => B_11_port);
   U69 : OAI21_X1 port map( B1 => n192, B2 => n63, A => n3, ZN => B_10_port);
   U70 : OAI21_X1 port map( B1 => n192, B2 => n39, A => n3, ZN => B_2_port);
   U71 : OAI21_X1 port map( B1 => n193, B2 => n116, A => n3, ZN => B_1_port);
   U72 : OAI221_X1 port map( B1 => n27, B2 => n11, C1 => n28, C2 => n191, A => 
                           n29, ZN => B_30_port);
   U73 : OAI221_X1 port map( B1 => n40, B2 => n11, C1 => n41, C2 => n191, A => 
                           n42, ZN => B_29_port);
   U74 : OAI221_X1 port map( B1 => n47, B2 => n11, C1 => n48, C2 => n191, A => 
                           n49, ZN => B_28_port);
   U75 : OAI221_X1 port map( B1 => n10, B2 => n55, C1 => n56, C2 => n191, A => 
                           n57, ZN => B_27_port);
   U76 : OAI221_X1 port map( B1 => n27, B2 => n55, C1 => n63, C2 => n191, A => 
                           n64, ZN => B_26_port);
   U77 : OAI221_X1 port map( B1 => n40, B2 => n55, C1 => n2, C2 => n191, A => 
                           n69, ZN => B_25_port);
   U78 : OAI221_X1 port map( B1 => n47, B2 => n55, C1 => n4, C2 => n191, A => 
                           n83, ZN => B_24_port);
   U79 : OAI221_X1 port map( B1 => n60, B2 => n55, C1 => n5, C2 => n191, A => 
                           n91, ZN => B_23_port);
   U80 : OAI221_X1 port map( B1 => n66, B2 => n55, C1 => n6, C2 => n191, A => 
                           n98, ZN => B_22_port);
   U81 : OAI221_X1 port map( B1 => n71, B2 => n55, C1 => n7, C2 => n191, A => 
                           n105, ZN => B_21_port);
   U82 : OAI221_X1 port map( B1 => n85, B2 => n55, C1 => n8, C2 => n191, A => 
                           n111, ZN => B_20_port);
   U83 : OAI221_X1 port map( B1 => n93, B2 => n55, C1 => n9, C2 => n191, A => 
                           n117, ZN => B_19_port);
   U84 : OAI221_X1 port map( B1 => n100, B2 => n55, C1 => n39, C2 => n191, A =>
                           n120, ZN => B_18_port);
   U85 : OAI221_X1 port map( B1 => n106, B2 => n55, C1 => n116, C2 => n191, A 
                           => n123, ZN => B_17_port);
   U86 : OAI221_X1 port map( B1 => n128, B2 => n11, C1 => n112, C2 => n55, A =>
                           n129, ZN => B_16_port);
   U87 : OAI21_X1 port map( B1 => n124, B2 => n188, A => n107, ZN => n113);
   U88 : AOI221_X1 port map( B1 => n14, B2 => n86, C1 => n18, C2 => n87, A => 
                           n130, ZN => n129);
   U89 : INV_X1 port map( A => n3, ZN => n130);
   U90 : NOR2_X1 port map( A1 => n188, A2 => n107, ZN => n80);
   U91 : NAND2_X1 port map( A1 => n186, A2 => n187, ZN => n34);
   U92 : AND2_X1 port map( A1 => n131, A2 => n188, ZN => n18);
   U93 : AND2_X1 port map( A1 => SH(3), A2 => n188, ZN => n78);
   U94 : AOI21_X1 port map( B1 => n86, B2 => n75, A => n113, ZN => n8);
   U95 : AOI21_X1 port map( B1 => n94, B2 => n75, A => n113, ZN => n9);
   U96 : AOI21_X1 port map( B1 => n101, B2 => n75, A => n113, ZN => n39);
   U97 : AOI21_X1 port map( B1 => n79, B2 => n75, A => n113, ZN => n116);
   U98 : INV_X1 port map( A => n107, ZN => n88);
   U99 : INV_X1 port map( A => n93, ZN => n15);
   U100 : INV_X1 port map( A => n100, ZN => n30);
   U101 : INV_X1 port map( A => n106, ZN => n43);
   U102 : INV_X1 port map( A => n112, ZN => n50);
   U103 : INV_X1 port map( A => n60, ZN => n19);
   U104 : INV_X1 port map( A => n66, ZN => n32);
   U105 : INV_X1 port map( A => n71, ZN => n45);
   U106 : INV_X1 port map( A => n85, ZN => n52);
   U107 : INV_X1 port map( A => n84, ZN => n128);
   U108 : AND2_X1 port map( A1 => SH(3), A2 => n191, ZN => n131);
   U109 : BUF_X1 port map( A => SH(4), Z => n190);
   U110 : BUF_X1 port map( A => SH(4), Z => n189);
   U111 : OAI221_X1 port map( B1 => n154, B2 => n20, C1 => n124, C2 => n22, A 
                           => n162, ZN => n94);
   U112 : AOI22_X1 port map( A1 => n25, A2 => A(2), B1 => A(3), B2 => n26, ZN 
                           => n162);
   U113 : OAI221_X1 port map( B1 => n33, B2 => n158, C1 => n34, C2 => n148, A 
                           => n159, ZN => n87);
   U114 : AOI22_X1 port map( A1 => A(6), A2 => n37, B1 => A(5), B2 => n38, ZN 
                           => n159);
   U115 : OAI221_X1 port map( B1 => n33, B2 => n165, C1 => n34, C2 => n158, A 
                           => n166, ZN => n95);
   U116 : AOI22_X1 port map( A1 => A(5), A2 => n37, B1 => A(4), B2 => n38, ZN 
                           => n166);
   U117 : OAI221_X1 port map( B1 => n33, B2 => n143, C1 => n34, C2 => n144, A 
                           => n145, ZN => n72);
   U118 : INV_X1 port map( A => A(4), ZN => n143);
   U119 : AOI22_X1 port map( A1 => A(3), A2 => n37, B1 => A(2), B2 => n38, ZN 
                           => n145);
   U120 : OAI221_X1 port map( B1 => n33, B2 => n156, C1 => n34, C2 => n146, A 
                           => n157, ZN => n84);
   U121 : AOI22_X1 port map( A1 => A(10), A2 => n37, B1 => A(9), B2 => n38, ZN 
                           => n157);
   U122 : OAI221_X1 port map( B1 => n33, B2 => n163, C1 => n34, C2 => n156, A 
                           => n164, ZN => n92);
   U123 : AOI22_X1 port map( A1 => A(9), A2 => n37, B1 => A(8), B2 => n38, ZN 
                           => n164);
   U124 : OAI221_X1 port map( B1 => n33, B2 => n149, C1 => n34, C2 => n163, A 
                           => n170, ZN => n99);
   U125 : AOI22_X1 port map( A1 => A(8), A2 => n37, B1 => A(7), B2 => n38, ZN 
                           => n170);
   U126 : OAI221_X1 port map( B1 => n33, B2 => n148, C1 => n34, C2 => n149, A 
                           => n150, ZN => n74);
   U127 : AOI22_X1 port map( A1 => A(7), A2 => n37, B1 => A(6), B2 => n38, ZN 
                           => n150);
   U128 : OAI221_X1 port map( B1 => n33, B2 => n127, C1 => n34, C2 => n122, A 
                           => n137, ZN => n59);
   U129 : AOI22_X1 port map( A1 => A(13), A2 => n37, B1 => A(12), B2 => n38, ZN
                           => n137);
   U130 : OAI221_X1 port map( B1 => n33, B2 => n133, C1 => n34, C2 => n127, A 
                           => n140, ZN => n65);
   U131 : AOI22_X1 port map( A1 => A(12), A2 => n37, B1 => A(11), B2 => n38, ZN
                           => n140);
   U132 : OAI221_X1 port map( B1 => n33, B2 => n146, C1 => n34, C2 => n133, A 
                           => n147, ZN => n70);
   U133 : AOI22_X1 port map( A1 => A(11), A2 => n37, B1 => A(10), B2 => n38, ZN
                           => n147);
   U134 : OAI221_X1 port map( B1 => n20, B2 => n153, C1 => n154, C2 => n22, A 
                           => n155, ZN => n86);
   U135 : AOI22_X1 port map( A1 => n25, A2 => A(3), B1 => A(4), B2 => n26, ZN 
                           => n155);
   U136 : AOI221_X1 port map( B1 => n25, B2 => A(26), C1 => n26, C2 => A(27), A
                           => n61, ZN => n10);
   U137 : INV_X1 port map( A => n62, ZN => n61);
   U138 : AOI22_X1 port map( A1 => A(25), A2 => n37, B1 => A(24), B2 => n38, ZN
                           => n62);
   U139 : AOI221_X1 port map( B1 => n25, B2 => A(25), C1 => n26, C2 => A(26), A
                           => n67, ZN => n27);
   U140 : INV_X1 port map( A => n68, ZN => n67);
   U141 : AOI22_X1 port map( A1 => A(24), A2 => n37, B1 => A(23), B2 => n38, ZN
                           => n68);
   U143 : AOI221_X1 port map( B1 => n25, B2 => A(24), C1 => n26, C2 => A(25), A
                           => n81, ZN => n40);
   U144 : INV_X1 port map( A => n82, ZN => n81);
   U145 : AOI22_X1 port map( A1 => A(23), A2 => n37, B1 => A(22), B2 => n38, ZN
                           => n82);
   U146 : AOI221_X1 port map( B1 => n25, B2 => A(23), C1 => n26, C2 => A(24), A
                           => n89, ZN => n47);
   U147 : INV_X1 port map( A => n90, ZN => n89);
   U148 : AOI22_X1 port map( A1 => A(22), A2 => n37, B1 => A(21), B2 => n38, ZN
                           => n90);
   U149 : AOI221_X1 port map( B1 => n25, B2 => A(22), C1 => n26, C2 => A(23), A
                           => n96, ZN => n60);
   U150 : INV_X1 port map( A => n97, ZN => n96);
   U151 : AOI22_X1 port map( A1 => A(21), A2 => n37, B1 => A(20), B2 => n38, ZN
                           => n97);
   U152 : AOI221_X1 port map( B1 => n25, B2 => A(21), C1 => n26, C2 => A(22), A
                           => n103, ZN => n66);
   U153 : INV_X1 port map( A => n104, ZN => n103);
   U154 : AOI22_X1 port map( A1 => A(20), A2 => n37, B1 => A(19), B2 => n38, ZN
                           => n104);
   U155 : AOI221_X1 port map( B1 => n25, B2 => A(20), C1 => n26, C2 => A(21), A
                           => n108, ZN => n71);
   U156 : OAI22_X1 port map( A1 => n109, A2 => n20, B1 => n110, B2 => n22, ZN 
                           => n108);
   U157 : INV_X1 port map( A => A(19), ZN => n109);
   U158 : AOI221_X1 port map( B1 => n25, B2 => A(19), C1 => n26, C2 => A(20), A
                           => n114, ZN => n85);
   U159 : OAI22_X1 port map( A1 => n110, A2 => n20, B1 => n115, B2 => n22, ZN 
                           => n114);
   U160 : AOI221_X1 port map( B1 => n25, B2 => A(18), C1 => n26, C2 => A(19), A
                           => n118, ZN => n93);
   U161 : OAI22_X1 port map( A1 => n115, A2 => n20, B1 => n119, B2 => n22, ZN 
                           => n118);
   U162 : AOI221_X1 port map( B1 => n25, B2 => A(17), C1 => n26, C2 => A(18), A
                           => n121, ZN => n100);
   U163 : OAI22_X1 port map( A1 => n119, A2 => n20, B1 => n122, B2 => n22, ZN 
                           => n121);
   U164 : AOI221_X1 port map( B1 => n25, B2 => A(16), C1 => n26, C2 => A(17), A
                           => n126, ZN => n106);
   U165 : OAI22_X1 port map( A1 => n122, A2 => n20, B1 => n127, B2 => n22, ZN 
                           => n126);
   U166 : AOI221_X1 port map( B1 => n25, B2 => A(15), C1 => n26, C2 => A(16), A
                           => n132, ZN => n112);
   U167 : OAI22_X1 port map( A1 => n127, A2 => n20, B1 => n133, B2 => n22, ZN 
                           => n132);
   U168 : AOI222_X1 port map( A1 => n14, A2 => n15, B1 => n16, B2 => n17, C1 =>
                           n18, C2 => n19, ZN => n13);
   U169 : OAI221_X1 port map( B1 => n20, B2 => n21, C1 => n22, C2 => n23, A => 
                           n24, ZN => n17);
   U170 : AOI22_X1 port map( A1 => A(30), A2 => n25, B1 => A(31), B2 => n26, ZN
                           => n24);
   U171 : AOI222_X1 port map( A1 => n14, A2 => n30, B1 => n16, B2 => n31, C1 =>
                           n18, C2 => n32, ZN => n29);
   U172 : OAI221_X1 port map( B1 => n33, B2 => n21, C1 => n34, C2 => n35, A => 
                           n36, ZN => n31);
   U173 : INV_X1 port map( A => A(30), ZN => n35);
   U174 : AOI22_X1 port map( A1 => A(28), A2 => n37, B1 => A(27), B2 => n38, ZN
                           => n36);
   U175 : AOI222_X1 port map( A1 => n14, A2 => n43, B1 => n16, B2 => n44, C1 =>
                           n18, C2 => n45, ZN => n42);
   U176 : OAI221_X1 port map( B1 => n33, B2 => n23, C1 => n34, C2 => n21, A => 
                           n46, ZN => n44);
   U177 : AOI22_X1 port map( A1 => A(27), A2 => n37, B1 => A(26), B2 => n38, ZN
                           => n46);
   U178 : AOI222_X1 port map( A1 => n14, A2 => n50, B1 => n16, B2 => n51, C1 =>
                           n18, C2 => n52, ZN => n49);
   U179 : OAI221_X1 port map( B1 => n33, B2 => n53, C1 => n34, C2 => n23, A => 
                           n54, ZN => n51);
   U180 : INV_X1 port map( A => A(27), ZN => n53);
   U181 : AOI22_X1 port map( A1 => A(26), A2 => n37, B1 => A(25), B2 => n38, ZN
                           => n54);
   U182 : NAND2_X1 port map( A1 => SH(1), A2 => n186, ZN => n20);
   U183 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n22);
   U184 : AND2_X1 port map( A1 => n131, A2 => SH(2), ZN => n14);
   U185 : NAND2_X1 port map( A1 => SH(3), A2 => A(0), ZN => n107);
   U186 : INV_X1 port map( A => n171, ZN => n102);
   U187 : AOI221_X1 port map( B1 => n37, B2 => A(4), C1 => A(3), C2 => n38, A 
                           => n172, ZN => n171);
   U188 : OAI22_X1 port map( A1 => n144, A2 => n33, B1 => n165, B2 => n34, ZN 
                           => n172);
   U189 : INV_X1 port map( A => A(14), ZN => n127);
   U190 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n136);
   U191 : INV_X1 port map( A => A(1), ZN => n154);
   U192 : INV_X1 port map( A => A(28), ZN => n23);
   U193 : INV_X1 port map( A => A(15), ZN => n122);
   U194 : INV_X1 port map( A => A(13), ZN => n133);
   U195 : INV_X1 port map( A => A(29), ZN => n21);
   U196 : INV_X1 port map( A => A(0), ZN => n124);
   U197 : INV_X1 port map( A => A(5), ZN => n144);
   U198 : INV_X1 port map( A => A(10), ZN => n163);
   U199 : INV_X1 port map( A => A(9), ZN => n149);
   U200 : INV_X1 port map( A => A(8), ZN => n148);
   U201 : INV_X1 port map( A => A(7), ZN => n158);
   U202 : INV_X1 port map( A => A(12), ZN => n146);
   U203 : INV_X1 port map( A => A(11), ZN => n156);
   U204 : INV_X1 port map( A => A(18), ZN => n110);
   U205 : INV_X1 port map( A => A(17), ZN => n115);
   U206 : INV_X1 port map( A => A(16), ZN => n119);
   U207 : INV_X1 port map( A => A(6), ZN => n165);
   U208 : INV_X1 port map( A => A(2), ZN => n153);
   U209 : INV_X1 port map( A => SH(0), ZN => n186);
   U210 : INV_X1 port map( A => SH(1), ZN => n187);
   U211 : INV_X1 port map( A => SH(2), ZN => n188);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Shifter_NBIT32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end Shifter_NBIT32_DW01_ash_0;

architecture SYN_mx2 of Shifter_NBIT32_DW01_ash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n3, n4, n5, n6, n7, n8, n9, n10, n28, n29, n30, n31, n32
      , n33, n34 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => SH(4), Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n33, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n33, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n33, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n33, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => SH(4), Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n33, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n33, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => SH(4), Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n33, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => SH(4), Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n33, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => SH(4), Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n33, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => SH(4), Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => SH(4), Z => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n31, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n31, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n31, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n31, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n31, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n31, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n31, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n31, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n31, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n31, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n31, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n31, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n31, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => SH(3), Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n31, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n31, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => SH(3), Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n31, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n31, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n31, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n31, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n31, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => SH(2), Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => SH(2), Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => SH(2), Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => SH(2), Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => SH(2), Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => SH(2), Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => SH(2), Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           SH(2), Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           SH(2), Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           SH(2), Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           SH(2), Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => SH(1), Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => SH(1), Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => SH(1), Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => SH(1), Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           SH(1), Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           SH(1), Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           SH(1), Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           SH(1), Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           SH(1), Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           SH(1), Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           SH(1), Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           SH(1), Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => SH(0), Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => SH(0), Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => SH(0), Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => SH(0), Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => SH(0), Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => SH(0), Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => SH(0), Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => SH(0), Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => SH(0), Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => SH(0), Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => SH(0), Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => SH(0), Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => SH(0), Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => SH(0), Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => SH(0), Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => SH(0), Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => SH(0), Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => SH(0), Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => SH(0), Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => SH(0), Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => SH(0), Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => SH(0), Z => 
                           ML_int_1_1_port);
   U3 : INV_X1 port map( A => n3, ZN => ML_int_4_7_port);
   U4 : INV_X1 port map( A => n4, ZN => ML_int_4_6_port);
   U5 : INV_X1 port map( A => n5, ZN => ML_int_4_5_port);
   U6 : INV_X1 port map( A => n6, ZN => ML_int_4_4_port);
   U7 : INV_X1 port map( A => n7, ZN => ML_int_4_3_port);
   U8 : INV_X1 port map( A => n8, ZN => ML_int_4_2_port);
   U9 : INV_X1 port map( A => n9, ZN => ML_int_4_1_port);
   U10 : INV_X1 port map( A => n10, ZN => ML_int_4_0_port);
   U11 : INV_X1 port map( A => n34, ZN => n33);
   U12 : INV_X1 port map( A => n32, ZN => n31);
   U13 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n32, ZN => n10);
   U14 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n32, ZN => n3);
   U15 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n32, ZN => n4);
   U16 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n32, ZN => n5);
   U17 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n32, ZN => n6);
   U18 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n32, ZN => n7);
   U19 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n32, ZN => n8);
   U20 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n32, ZN => n9);
   U21 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n34, ZN => B(9));
   U22 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n34, ZN => B(8));
   U23 : NOR2_X1 port map( A1 => n33, A2 => n3, ZN => B(7));
   U24 : NOR2_X1 port map( A1 => n33, A2 => n4, ZN => B(6));
   U25 : NOR2_X1 port map( A1 => n33, A2 => n5, ZN => B(5));
   U26 : NOR2_X1 port map( A1 => n33, A2 => n6, ZN => B(4));
   U27 : NOR2_X1 port map( A1 => n33, A2 => n7, ZN => B(3));
   U28 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n34, ZN => B(15));
   U29 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n34, ZN => B(14));
   U30 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n34, ZN => B(13));
   U31 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n34, ZN => B(12));
   U32 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n34, ZN => B(11));
   U33 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n34, ZN => B(10));
   U34 : NOR2_X1 port map( A1 => n33, A2 => n8, ZN => B(2));
   U35 : NOR2_X1 port map( A1 => n33, A2 => n9, ZN => B(1));
   U36 : INV_X1 port map( A => SH(4), ZN => n34);
   U37 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n30, ZN => 
                           ML_int_3_3_port);
   U38 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n30, ZN => 
                           ML_int_3_2_port);
   U39 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n30, ZN => 
                           ML_int_3_0_port);
   U40 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n30, ZN => 
                           ML_int_3_1_port);
   U41 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n29, ZN => 
                           ML_int_2_0_port);
   U42 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n29, ZN => 
                           ML_int_2_1_port);
   U43 : NOR2_X1 port map( A1 => n33, A2 => n10, ZN => B(0));
   U44 : INV_X1 port map( A => SH(1), ZN => n29);
   U45 : INV_X1 port map( A => SH(0), ZN => n28);
   U46 : INV_X1 port map( A => SH(2), ZN => n30);
   U47 : AND2_X1 port map( A1 => A(0), A2 => n28, ZN => ML_int_1_0_port);
   U48 : INV_X1 port map( A => SH(3), ZN => n32);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity DIVIDER_N_op32_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end DIVIDER_N_op32_DW01_sub_0;

architecture SYN_rpl of DIVIDER_N_op32_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, DIFF_2_port, 
      DIFF_1_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, B_not_31_port, 
      B_not_30_port, B_not_29_port, B_not_28_port, B_not_27_port, B_not_26_port
      , B_not_25_port, B_not_24_port, B_not_23_port, B_not_22_port, 
      B_not_21_port, B_not_20_port, B_not_19_port, B_not_18_port, B_not_17_port
      , B_not_16_port, B_not_15_port, B_not_14_port, B_not_13_port, 
      B_not_12_port, B_not_11_port, B_not_10_port, B_not_9_port, B_not_8_port, 
      B_not_7_port, B_not_6_port, B_not_5_port, B_not_4_port, B_not_3_port, 
      B_not_2_port, B_not_1_port, net88787 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U2_31 : FA_X1 port map( A => A(31), B => B_not_31_port, CI => carry_31_port,
                           CO => net88787, S => DIFF_31_port);
   U2_30 : FA_X1 port map( A => A(30), B => B_not_30_port, CI => carry_30_port,
                           CO => carry_31_port, S => DIFF_30_port);
   U2_29 : FA_X1 port map( A => A(29), B => B_not_29_port, CI => carry_29_port,
                           CO => carry_30_port, S => DIFF_29_port);
   U2_28 : FA_X1 port map( A => A(28), B => B_not_28_port, CI => carry_28_port,
                           CO => carry_29_port, S => DIFF_28_port);
   U2_27 : FA_X1 port map( A => A(27), B => B_not_27_port, CI => carry_27_port,
                           CO => carry_28_port, S => DIFF_27_port);
   U2_26 : FA_X1 port map( A => A(26), B => B_not_26_port, CI => carry_26_port,
                           CO => carry_27_port, S => DIFF_26_port);
   U2_25 : FA_X1 port map( A => A(25), B => B_not_25_port, CI => carry_25_port,
                           CO => carry_26_port, S => DIFF_25_port);
   U2_24 : FA_X1 port map( A => A(24), B => B_not_24_port, CI => carry_24_port,
                           CO => carry_25_port, S => DIFF_24_port);
   U2_23 : FA_X1 port map( A => A(23), B => B_not_23_port, CI => carry_23_port,
                           CO => carry_24_port, S => DIFF_23_port);
   U2_22 : FA_X1 port map( A => A(22), B => B_not_22_port, CI => carry_22_port,
                           CO => carry_23_port, S => DIFF_22_port);
   U2_21 : FA_X1 port map( A => A(21), B => B_not_21_port, CI => carry_21_port,
                           CO => carry_22_port, S => DIFF_21_port);
   U2_20 : FA_X1 port map( A => A(20), B => B_not_20_port, CI => carry_20_port,
                           CO => carry_21_port, S => DIFF_20_port);
   U2_19 : FA_X1 port map( A => A(19), B => B_not_19_port, CI => carry_19_port,
                           CO => carry_20_port, S => DIFF_19_port);
   U2_18 : FA_X1 port map( A => A(18), B => B_not_18_port, CI => carry_18_port,
                           CO => carry_19_port, S => DIFF_18_port);
   U2_17 : FA_X1 port map( A => A(17), B => B_not_17_port, CI => carry_17_port,
                           CO => carry_18_port, S => DIFF_17_port);
   U2_16 : FA_X1 port map( A => A(16), B => B_not_16_port, CI => carry_16_port,
                           CO => carry_17_port, S => DIFF_16_port);
   U2_15 : FA_X1 port map( A => A(15), B => B_not_15_port, CI => carry_15_port,
                           CO => carry_16_port, S => DIFF_15_port);
   U2_14 : FA_X1 port map( A => A(14), B => B_not_14_port, CI => carry_14_port,
                           CO => carry_15_port, S => DIFF_14_port);
   U2_13 : FA_X1 port map( A => A(13), B => B_not_13_port, CI => carry_13_port,
                           CO => carry_14_port, S => DIFF_13_port);
   U2_12 : FA_X1 port map( A => A(12), B => B_not_12_port, CI => carry_12_port,
                           CO => carry_13_port, S => DIFF_12_port);
   U2_11 : FA_X1 port map( A => A(11), B => B_not_11_port, CI => carry_11_port,
                           CO => carry_12_port, S => DIFF_11_port);
   U2_10 : FA_X1 port map( A => A(10), B => B_not_10_port, CI => carry_10_port,
                           CO => carry_11_port, S => DIFF_10_port);
   U2_9 : FA_X1 port map( A => A(9), B => B_not_9_port, CI => carry_9_port, CO 
                           => carry_10_port, S => DIFF_9_port);
   U2_8 : FA_X1 port map( A => A(8), B => B_not_8_port, CI => carry_8_port, CO 
                           => carry_9_port, S => DIFF_8_port);
   U2_7 : FA_X1 port map( A => A(7), B => B_not_7_port, CI => carry_7_port, CO 
                           => carry_8_port, S => DIFF_7_port);
   U2_6 : FA_X1 port map( A => A(6), B => B_not_6_port, CI => carry_6_port, CO 
                           => carry_7_port, S => DIFF_6_port);
   U2_5 : FA_X1 port map( A => A(5), B => B_not_5_port, CI => carry_5_port, CO 
                           => carry_6_port, S => DIFF_5_port);
   U2_4 : FA_X1 port map( A => A(4), B => B_not_4_port, CI => carry_4_port, CO 
                           => carry_5_port, S => DIFF_4_port);
   U2_3 : FA_X1 port map( A => A(3), B => B_not_3_port, CI => carry_3_port, CO 
                           => carry_4_port, S => DIFF_3_port);
   U2_2 : FA_X1 port map( A => A(2), B => B_not_2_port, CI => carry_2_port, CO 
                           => carry_3_port, S => DIFF_2_port);
   U2_1 : FA_X1 port map( A => A(1), B => B_not_1_port, CI => carry_1_port, CO 
                           => carry_2_port, S => DIFF_1_port);
   U1 : INV_X1 port map( A => B(0), ZN => carry_1_port);
   U2 : INV_X1 port map( A => B(1), ZN => B_not_1_port);
   U3 : INV_X1 port map( A => B(2), ZN => B_not_2_port);
   U4 : INV_X1 port map( A => B(3), ZN => B_not_3_port);
   U5 : INV_X1 port map( A => B(4), ZN => B_not_4_port);
   U6 : INV_X1 port map( A => B(5), ZN => B_not_5_port);
   U7 : INV_X1 port map( A => B(6), ZN => B_not_6_port);
   U8 : INV_X1 port map( A => B(7), ZN => B_not_7_port);
   U9 : INV_X1 port map( A => B(8), ZN => B_not_8_port);
   U10 : INV_X1 port map( A => B(9), ZN => B_not_9_port);
   U11 : INV_X1 port map( A => B(10), ZN => B_not_10_port);
   U12 : INV_X1 port map( A => B(11), ZN => B_not_11_port);
   U13 : INV_X1 port map( A => B(12), ZN => B_not_12_port);
   U14 : INV_X1 port map( A => B(13), ZN => B_not_13_port);
   U15 : INV_X1 port map( A => B(14), ZN => B_not_14_port);
   U16 : INV_X1 port map( A => B(15), ZN => B_not_15_port);
   U17 : INV_X1 port map( A => B(16), ZN => B_not_16_port);
   U18 : INV_X1 port map( A => B(17), ZN => B_not_17_port);
   U19 : INV_X1 port map( A => B(18), ZN => B_not_18_port);
   U20 : INV_X1 port map( A => B(19), ZN => B_not_19_port);
   U21 : INV_X1 port map( A => B(20), ZN => B_not_20_port);
   U22 : INV_X1 port map( A => B(21), ZN => B_not_21_port);
   U23 : INV_X1 port map( A => B(22), ZN => B_not_22_port);
   U24 : INV_X1 port map( A => B(23), ZN => B_not_23_port);
   U25 : INV_X1 port map( A => B(24), ZN => B_not_24_port);
   U26 : INV_X1 port map( A => B(25), ZN => B_not_25_port);
   U27 : INV_X1 port map( A => B(26), ZN => B_not_26_port);
   U28 : INV_X1 port map( A => B(27), ZN => B_not_27_port);
   U29 : INV_X1 port map( A => B(28), ZN => B_not_28_port);
   U30 : INV_X1 port map( A => B(29), ZN => B_not_29_port);
   U31 : INV_X1 port map( A => B(30), ZN => B_not_30_port);
   U32 : INV_X1 port map( A => B(31), ZN => B_not_31_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity DIVIDER_N_op32_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end DIVIDER_N_op32_DW01_inc_0;

architecture SYN_rpl of DIVIDER_N_op32_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity cu_lower_mux is

   port( EX_MEM_write, MEM_WB_write : in std_logic;  EX_MEM_Rd, ID_EX_Rt, 
         MEM_WB_Rd : in std_logic_vector (4 downto 0);  sel_lower_mux : out 
         std_logic_vector (1 downto 0));

end cu_lower_mux;

architecture SYN_Behavioral of cu_lower_mux is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14 : std_logic;

begin
   
   U11 : XOR2_X1 port map( A => MEM_WB_Rd(1), B => ID_EX_Rt(1), Z => n5);
   U12 : XOR2_X1 port map( A => MEM_WB_Rd(2), B => ID_EX_Rt(2), Z => n4);
   U13 : XOR2_X1 port map( A => MEM_WB_Rd(3), B => ID_EX_Rt(3), Z => n3);
   U14 : XOR2_X1 port map( A => ID_EX_Rt(3), B => EX_MEM_Rd(3), Z => n14);
   U15 : XOR2_X1 port map( A => ID_EX_Rt(2), B => EX_MEM_Rd(2), Z => n13);
   U16 : XOR2_X1 port map( A => ID_EX_Rt(4), B => EX_MEM_Rd(4), Z => n12);
   U2 : INV_X1 port map( A => n8, ZN => sel_lower_mux(0));
   U3 : NOR4_X1 port map( A1 => n2, A2 => n3, A3 => n4, A4 => n5, ZN => 
                           sel_lower_mux(1));
   U4 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => MEM_WB_write, A4 => n8, ZN
                           => n2);
   U5 : NAND4_X1 port map( A1 => n9, A2 => EX_MEM_write, A3 => n10, A4 => n11, 
                           ZN => n8);
   U6 : XNOR2_X1 port map( A => ID_EX_Rt(1), B => EX_MEM_Rd(1), ZN => n9);
   U7 : XNOR2_X1 port map( A => ID_EX_Rt(0), B => EX_MEM_Rd(0), ZN => n10);
   U8 : NOR3_X1 port map( A1 => n12, A2 => n13, A3 => n14, ZN => n11);
   U9 : XNOR2_X1 port map( A => ID_EX_Rt(0), B => MEM_WB_Rd(0), ZN => n7);
   U10 : XNOR2_X1 port map( A => ID_EX_Rt(4), B => MEM_WB_Rd(4), ZN => n6);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity cu_upper_mux is

   port( EX_MEM_write, MEM_WB_write : in std_logic;  MEM_WB_Rd, EX_MEM_Rd, 
         ID_EX_Rs : in std_logic_vector (4 downto 0);  sel_upper_mux : out 
         std_logic_vector (1 downto 0));

end cu_upper_mux;

architecture SYN_Behavioral of cu_upper_mux is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14 : std_logic;

begin
   
   U11 : XOR2_X1 port map( A => MEM_WB_Rd(1), B => ID_EX_Rs(1), Z => n5);
   U12 : XOR2_X1 port map( A => MEM_WB_Rd(2), B => ID_EX_Rs(2), Z => n4);
   U13 : XOR2_X1 port map( A => MEM_WB_Rd(3), B => ID_EX_Rs(3), Z => n3);
   U14 : XOR2_X1 port map( A => ID_EX_Rs(3), B => EX_MEM_Rd(3), Z => n14);
   U15 : XOR2_X1 port map( A => ID_EX_Rs(2), B => EX_MEM_Rd(2), Z => n13);
   U16 : XOR2_X1 port map( A => ID_EX_Rs(4), B => EX_MEM_Rd(4), Z => n12);
   U2 : INV_X1 port map( A => n8, ZN => sel_upper_mux(0));
   U3 : NOR4_X1 port map( A1 => n2, A2 => n3, A3 => n4, A4 => n5, ZN => 
                           sel_upper_mux(1));
   U4 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => MEM_WB_write, A4 => n8, ZN
                           => n2);
   U5 : NAND4_X1 port map( A1 => n9, A2 => EX_MEM_write, A3 => n10, A4 => n11, 
                           ZN => n8);
   U6 : XNOR2_X1 port map( A => ID_EX_Rs(1), B => EX_MEM_Rd(1), ZN => n9);
   U7 : XNOR2_X1 port map( A => ID_EX_Rs(0), B => EX_MEM_Rd(0), ZN => n10);
   U8 : NOR3_X1 port map( A1 => n12, A2 => n13, A3 => n14, ZN => n11);
   U9 : XNOR2_X1 port map( A => ID_EX_Rs(0), B => MEM_WB_Rd(0), ZN => n7);
   U10 : XNOR2_X1 port map( A => ID_EX_Rs(4), B => MEM_WB_Rd(4), ZN => n6);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Adder is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  O : out
         std_logic_vector (31 downto 0);  CO : out std_logic);

end Adder;

architecture SYN_Behavioral of Adder is

   component Adder_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal CO_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, O_0_port, 
      net166339 : std_logic;

begin
   O <= ( CO_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, O_0_port );
   CO <= CO_port;
   
   add_1_root_add_24_2 : Adder_DW01_add_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => CI, SUM(31) => CO_port,
                           SUM(30) => O_30_port, SUM(29) => O_29_port, SUM(28) 
                           => O_28_port, SUM(27) => O_27_port, SUM(26) => 
                           O_26_port, SUM(25) => O_25_port, SUM(24) => 
                           O_24_port, SUM(23) => O_23_port, SUM(22) => 
                           O_22_port, SUM(21) => O_21_port, SUM(20) => 
                           O_20_port, SUM(19) => O_19_port, SUM(18) => 
                           O_18_port, SUM(17) => O_17_port, SUM(16) => 
                           O_16_port, SUM(15) => O_15_port, SUM(14) => 
                           O_14_port, SUM(13) => O_13_port, SUM(12) => 
                           O_12_port, SUM(11) => O_11_port, SUM(10) => 
                           O_10_port, SUM(9) => O_9_port, SUM(8) => O_8_port, 
                           SUM(7) => O_7_port, SUM(6) => O_6_port, SUM(5) => 
                           O_5_port, SUM(4) => O_4_port, SUM(3) => O_3_port, 
                           SUM(2) => O_2_port, SUM(1) => O_1_port, SUM(0) => 
                           O_0_port, CO => net166339);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity InstructionRegister is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end InstructionRegister;

architecture SYN_Behavioral of InstructionRegister is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n37, n39, n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n31, n32, n33, n34, n35, n38, n40, n42, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191 : std_logic;

begin
   
   R_reg_31_inst : DFF_X1 port map( D => n100, CK => n191, Q => o(31), QN => 
                           n37);
   R_reg_30_inst : DFF_X1 port map( D => n99, CK => n191, Q => o(30), QN => n33
                           );
   R_reg_29_inst : DFF_X1 port map( D => n98, CK => n191, Q => o(29), QN => n39
                           );
   R_reg_28_inst : DFF_X1 port map( D => n97, CK => n191, Q => o(28), QN => n32
                           );
   R_reg_27_inst : DFF_X1 port map( D => n96, CK => n191, Q => o(27), QN => n41
                           );
   R_reg_26_inst : DFF_X1 port map( D => n95, CK => n191, Q => o(26), QN => n31
                           );
   R_reg_25_inst : DFF_X1 port map( D => n94, CK => n189, Q => o(25), QN => n43
                           );
   R_reg_24_inst : DFF_X1 port map( D => n93, CK => n191, Q => o(24), QN => n44
                           );
   R_reg_23_inst : DFF_X1 port map( D => n92, CK => n191, Q => o(23), QN => n45
                           );
   R_reg_22_inst : DFF_X1 port map( D => n91, CK => n191, Q => o(22), QN => n46
                           );
   R_reg_21_inst : DFF_X1 port map( D => n90, CK => n191, Q => o(21), QN => n47
                           );
   R_reg_20_inst : DFF_X1 port map( D => n89, CK => n190, Q => o(20), QN => n48
                           );
   R_reg_19_inst : DFF_X1 port map( D => n88, CK => n190, Q => o(19), QN => n49
                           );
   R_reg_18_inst : DFF_X1 port map( D => n87, CK => n190, Q => o(18), QN => n50
                           );
   R_reg_17_inst : DFF_X1 port map( D => n86, CK => n190, Q => o(17), QN => n51
                           );
   R_reg_16_inst : DFF_X1 port map( D => n85, CK => n190, Q => o(16), QN => n52
                           );
   R_reg_15_inst : DFF_X1 port map( D => n84, CK => n190, Q => o(15), QN => n53
                           );
   R_reg_14_inst : DFF_X1 port map( D => n83, CK => n190, Q => o(14), QN => n54
                           );
   R_reg_13_inst : DFF_X1 port map( D => n82, CK => n190, Q => o(13), QN => n55
                           );
   R_reg_12_inst : DFF_X1 port map( D => n81, CK => n190, Q => o(12), QN => n56
                           );
   R_reg_11_inst : DFF_X1 port map( D => n80, CK => n190, Q => o(11), QN => n57
                           );
   R_reg_10_inst : DFF_X1 port map( D => n79, CK => n190, Q => o(10), QN => n58
                           );
   R_reg_9_inst : DFF_X1 port map( D => n78, CK => n189, Q => o(9), QN => n59);
   R_reg_8_inst : DFF_X1 port map( D => n77, CK => n189, Q => o(8), QN => n60);
   R_reg_7_inst : DFF_X1 port map( D => n76, CK => n189, Q => o(7), QN => n61);
   R_reg_6_inst : DFF_X1 port map( D => n75, CK => n189, Q => o(6), QN => n62);
   R_reg_5_inst : DFF_X1 port map( D => n74, CK => n189, Q => o(5), QN => n63);
   R_reg_4_inst : DFF_X1 port map( D => n73, CK => n189, Q => o(4), QN => n64);
   R_reg_3_inst : DFF_X1 port map( D => n72, CK => n189, Q => o(3), QN => n65);
   R_reg_2_inst : DFF_X1 port map( D => n71, CK => n189, Q => o(2), QN => n66);
   R_reg_1_inst : DFF_X1 port map( D => n70, CK => n189, Q => o(1), QN => n67);
   R_reg_0_inst : DFF_X1 port map( D => n69, CK => n189, Q => o(0), QN => n68);
   U3 : BUF_X1 port map( A => n38, Z => n183);
   U4 : BUF_X1 port map( A => n38, Z => n182);
   U5 : BUF_X1 port map( A => n38, Z => n184);
   U6 : BUF_X1 port map( A => n34, Z => n185);
   U7 : BUF_X1 port map( A => n34, Z => n186);
   U8 : BUF_X1 port map( A => n34, Z => n187);
   U9 : NAND2_X1 port map( A1 => n188, A2 => n185, ZN => n38);
   U10 : BUF_X1 port map( A => clock, Z => n190);
   U11 : BUF_X1 port map( A => clock, Z => n189);
   U12 : BUF_X1 port map( A => clock, Z => n191);
   U13 : OAI22_X1 port map( A1 => n187, A2 => n68, B1 => n184, B2 => n128, ZN 
                           => n69);
   U14 : INV_X1 port map( A => i(0), ZN => n128);
   U15 : OAI22_X1 port map( A1 => n187, A2 => n67, B1 => n184, B2 => n127, ZN 
                           => n70);
   U16 : INV_X1 port map( A => i(1), ZN => n127);
   U17 : OAI22_X1 port map( A1 => n187, A2 => n66, B1 => n184, B2 => n126, ZN 
                           => n71);
   U18 : INV_X1 port map( A => i(2), ZN => n126);
   U19 : OAI22_X1 port map( A1 => n187, A2 => n65, B1 => n184, B2 => n125, ZN 
                           => n72);
   U20 : INV_X1 port map( A => i(3), ZN => n125);
   U21 : OAI22_X1 port map( A1 => n187, A2 => n64, B1 => n183, B2 => n124, ZN 
                           => n73);
   U22 : INV_X1 port map( A => i(4), ZN => n124);
   U23 : OAI22_X1 port map( A1 => n187, A2 => n63, B1 => n183, B2 => n123, ZN 
                           => n74);
   U24 : INV_X1 port map( A => i(5), ZN => n123);
   U25 : OAI22_X1 port map( A1 => n187, A2 => n62, B1 => n183, B2 => n122, ZN 
                           => n75);
   U26 : INV_X1 port map( A => i(6), ZN => n122);
   U27 : OAI22_X1 port map( A1 => n186, A2 => n61, B1 => n183, B2 => n121, ZN 
                           => n76);
   U28 : INV_X1 port map( A => i(7), ZN => n121);
   U29 : OAI22_X1 port map( A1 => n186, A2 => n60, B1 => n183, B2 => n120, ZN 
                           => n77);
   U30 : INV_X1 port map( A => i(8), ZN => n120);
   U31 : OAI22_X1 port map( A1 => n186, A2 => n59, B1 => n183, B2 => n119, ZN 
                           => n78);
   U32 : INV_X1 port map( A => i(9), ZN => n119);
   U33 : OAI22_X1 port map( A1 => n186, A2 => n58, B1 => n183, B2 => n118, ZN 
                           => n79);
   U34 : INV_X1 port map( A => i(10), ZN => n118);
   U35 : OAI22_X1 port map( A1 => n186, A2 => n57, B1 => n183, B2 => n117, ZN 
                           => n80);
   U36 : INV_X1 port map( A => i(11), ZN => n117);
   U37 : OAI22_X1 port map( A1 => n186, A2 => n56, B1 => n183, B2 => n116, ZN 
                           => n81);
   U38 : INV_X1 port map( A => i(12), ZN => n116);
   U39 : OAI22_X1 port map( A1 => n186, A2 => n55, B1 => n183, B2 => n115, ZN 
                           => n82);
   U40 : INV_X1 port map( A => i(13), ZN => n115);
   U41 : OAI22_X1 port map( A1 => n186, A2 => n54, B1 => n183, B2 => n114, ZN 
                           => n83);
   U42 : INV_X1 port map( A => i(14), ZN => n114);
   U43 : OAI22_X1 port map( A1 => n186, A2 => n53, B1 => n183, B2 => n113, ZN 
                           => n84);
   U44 : INV_X1 port map( A => i(15), ZN => n113);
   U45 : OAI22_X1 port map( A1 => n186, A2 => n52, B1 => n182, B2 => n112, ZN 
                           => n85);
   U46 : INV_X1 port map( A => i(16), ZN => n112);
   U47 : OAI22_X1 port map( A1 => n186, A2 => n51, B1 => n182, B2 => n111, ZN 
                           => n86);
   U48 : INV_X1 port map( A => i(17), ZN => n111);
   U49 : OAI22_X1 port map( A1 => n186, A2 => n50, B1 => n182, B2 => n110, ZN 
                           => n87);
   U50 : INV_X1 port map( A => i(18), ZN => n110);
   U51 : OAI22_X1 port map( A1 => n185, A2 => n49, B1 => n182, B2 => n109, ZN 
                           => n88);
   U52 : INV_X1 port map( A => i(19), ZN => n109);
   U53 : OAI22_X1 port map( A1 => n185, A2 => n48, B1 => n182, B2 => n108, ZN 
                           => n89);
   U54 : INV_X1 port map( A => i(20), ZN => n108);
   U55 : OAI22_X1 port map( A1 => n185, A2 => n47, B1 => n182, B2 => n107, ZN 
                           => n90);
   U56 : INV_X1 port map( A => i(21), ZN => n107);
   U57 : OAI22_X1 port map( A1 => n185, A2 => n46, B1 => n182, B2 => n106, ZN 
                           => n91);
   U58 : INV_X1 port map( A => i(22), ZN => n106);
   U59 : OAI22_X1 port map( A1 => n185, A2 => n45, B1 => n182, B2 => n105, ZN 
                           => n92);
   U60 : INV_X1 port map( A => i(23), ZN => n105);
   U61 : OAI22_X1 port map( A1 => n185, A2 => n44, B1 => n182, B2 => n104, ZN 
                           => n93);
   U62 : INV_X1 port map( A => i(24), ZN => n104);
   U63 : OAI22_X1 port map( A1 => n186, A2 => n43, B1 => n182, B2 => n103, ZN 
                           => n94);
   U64 : INV_X1 port map( A => i(25), ZN => n103);
   U65 : OAI22_X1 port map( A1 => n185, A2 => n41, B1 => n182, B2 => n101, ZN 
                           => n96);
   U66 : INV_X1 port map( A => i(27), ZN => n101);
   U67 : OAI22_X1 port map( A1 => n185, A2 => n39, B1 => n182, B2 => n40, ZN =>
                           n98);
   U68 : INV_X1 port map( A => i(29), ZN => n40);
   U69 : OAI22_X1 port map( A1 => n185, A2 => n37, B1 => n184, B2 => n129, ZN 
                           => n100);
   U70 : INV_X1 port map( A => i(31), ZN => n129);
   U71 : OAI211_X1 port map( C1 => n187, C2 => n31, A => n102, B => n188, ZN =>
                           n95);
   U72 : NAND2_X1 port map( A1 => i(26), A2 => n185, ZN => n102);
   U73 : OAI211_X1 port map( C1 => n187, C2 => n32, A => n42, B => n188, ZN => 
                           n97);
   U74 : NAND2_X1 port map( A1 => i(28), A2 => n185, ZN => n42);
   U75 : OAI211_X1 port map( C1 => n187, C2 => n33, A => n35, B => n188, ZN => 
                           n99);
   U76 : NAND2_X1 port map( A1 => i(30), A2 => n185, ZN => n35);
   U77 : OR2_X1 port map( A1 => reset, A2 => load, ZN => n34);
   U78 : INV_X1 port map( A => reset, ZN => n188);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity regWithLoad32bit is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end regWithLoad32bit;

architecture SYN_Behavioral of regWithLoad32bit is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n34, n35, n36, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196 : std_logic;

begin
   
   R_reg_31_inst : DFF_X1 port map( D => n100, CK => n194, Q => o(31), QN => 
                           n37);
   R_reg_30_inst : DFF_X1 port map( D => n99, CK => n194, Q => o(30), QN => n38
                           );
   R_reg_29_inst : DFF_X1 port map( D => n98, CK => n194, Q => o(29), QN => n39
                           );
   R_reg_28_inst : DFF_X1 port map( D => n97, CK => n194, Q => o(28), QN => n40
                           );
   R_reg_27_inst : DFF_X1 port map( D => n96, CK => n194, Q => o(27), QN => n41
                           );
   R_reg_26_inst : DFF_X1 port map( D => n95, CK => n194, Q => o(26), QN => n42
                           );
   R_reg_25_inst : DFF_X1 port map( D => n94, CK => n194, Q => o(25), QN => n43
                           );
   R_reg_24_inst : DFF_X1 port map( D => n93, CK => n194, Q => o(24), QN => n44
                           );
   R_reg_23_inst : DFF_X1 port map( D => n92, CK => n194, Q => o(23), QN => n45
                           );
   R_reg_22_inst : DFF_X1 port map( D => n91, CK => n194, Q => o(22), QN => n46
                           );
   R_reg_21_inst : DFF_X1 port map( D => n90, CK => n194, Q => o(21), QN => n47
                           );
   R_reg_20_inst : DFF_X1 port map( D => n89, CK => n195, Q => o(20), QN => n48
                           );
   R_reg_19_inst : DFF_X1 port map( D => n88, CK => n195, Q => o(19), QN => n49
                           );
   R_reg_18_inst : DFF_X1 port map( D => n87, CK => n195, Q => o(18), QN => n50
                           );
   R_reg_17_inst : DFF_X1 port map( D => n86, CK => n195, Q => o(17), QN => n51
                           );
   R_reg_16_inst : DFF_X1 port map( D => n85, CK => n195, Q => o(16), QN => n52
                           );
   R_reg_15_inst : DFF_X1 port map( D => n84, CK => n195, Q => o(15), QN => n53
                           );
   R_reg_14_inst : DFF_X1 port map( D => n83, CK => n195, Q => o(14), QN => n54
                           );
   R_reg_13_inst : DFF_X1 port map( D => n82, CK => n195, Q => o(13), QN => n55
                           );
   R_reg_12_inst : DFF_X1 port map( D => n81, CK => n195, Q => o(12), QN => n56
                           );
   R_reg_11_inst : DFF_X1 port map( D => n80, CK => n195, Q => o(11), QN => n57
                           );
   R_reg_10_inst : DFF_X1 port map( D => n79, CK => n195, Q => o(10), QN => n58
                           );
   R_reg_9_inst : DFF_X1 port map( D => n78, CK => n196, Q => o(9), QN => n59);
   R_reg_8_inst : DFF_X1 port map( D => n77, CK => n196, Q => o(8), QN => n60);
   R_reg_7_inst : DFF_X1 port map( D => n76, CK => n196, Q => o(7), QN => n61);
   R_reg_6_inst : DFF_X1 port map( D => n75, CK => n196, Q => o(6), QN => n62);
   R_reg_5_inst : DFF_X1 port map( D => n74, CK => n196, Q => o(5), QN => n63);
   R_reg_4_inst : DFF_X1 port map( D => n73, CK => n196, Q => o(4), QN => n64);
   R_reg_3_inst : DFF_X1 port map( D => n72, CK => n196, Q => o(3), QN => n65);
   R_reg_2_inst : DFF_X1 port map( D => n71, CK => n196, Q => o(2), QN => n66);
   R_reg_1_inst : DFF_X1 port map( D => n70, CK => n196, Q => o(1), QN => n67);
   R_reg_0_inst : DFF_X1 port map( D => n69, CK => n196, Q => o(0), QN => n68);
   U3 : BUF_X1 port map( A => n34, Z => n190);
   U4 : BUF_X1 port map( A => n34, Z => n191);
   U5 : BUF_X1 port map( A => n35, Z => n188);
   U6 : BUF_X1 port map( A => n35, Z => n187);
   U7 : BUF_X1 port map( A => n35, Z => n189);
   U8 : BUF_X1 port map( A => n34, Z => n192);
   U9 : BUF_X1 port map( A => clock, Z => n195);
   U10 : BUF_X1 port map( A => clock, Z => n194);
   U11 : BUF_X1 port map( A => clock, Z => n196);
   U12 : OAI22_X1 port map( A1 => n191, A2 => n45, B1 => n189, B2 => n107, ZN 
                           => n92);
   U13 : INV_X1 port map( A => i(23), ZN => n107);
   U14 : OAI22_X1 port map( A1 => n192, A2 => n44, B1 => n189, B2 => n106, ZN 
                           => n93);
   U15 : INV_X1 port map( A => i(24), ZN => n106);
   U16 : OAI22_X1 port map( A1 => n192, A2 => n43, B1 => n189, B2 => n105, ZN 
                           => n94);
   U17 : INV_X1 port map( A => i(25), ZN => n105);
   U18 : OAI22_X1 port map( A1 => n192, A2 => n42, B1 => n189, B2 => n104, ZN 
                           => n95);
   U19 : INV_X1 port map( A => i(26), ZN => n104);
   U20 : OAI22_X1 port map( A1 => n192, A2 => n41, B1 => n189, B2 => n103, ZN 
                           => n96);
   U21 : INV_X1 port map( A => i(27), ZN => n103);
   U22 : OAI22_X1 port map( A1 => n192, A2 => n40, B1 => n189, B2 => n102, ZN 
                           => n97);
   U23 : INV_X1 port map( A => i(28), ZN => n102);
   U24 : OAI22_X1 port map( A1 => n192, A2 => n39, B1 => n189, B2 => n101, ZN 
                           => n98);
   U25 : INV_X1 port map( A => i(29), ZN => n101);
   U26 : OAI22_X1 port map( A1 => n192, A2 => n38, B1 => n189, B2 => n36, ZN =>
                           n99);
   U27 : INV_X1 port map( A => i(30), ZN => n36);
   U28 : OAI22_X1 port map( A1 => n190, A2 => n68, B1 => n187, B2 => n130, ZN 
                           => n69);
   U29 : INV_X1 port map( A => i(0), ZN => n130);
   U30 : OAI22_X1 port map( A1 => n190, A2 => n67, B1 => n187, B2 => n129, ZN 
                           => n70);
   U31 : INV_X1 port map( A => i(1), ZN => n129);
   U32 : OAI22_X1 port map( A1 => n190, A2 => n66, B1 => n187, B2 => n128, ZN 
                           => n71);
   U33 : INV_X1 port map( A => i(2), ZN => n128);
   U34 : OAI22_X1 port map( A1 => n190, A2 => n65, B1 => n187, B2 => n127, ZN 
                           => n72);
   U35 : INV_X1 port map( A => i(3), ZN => n127);
   U36 : OAI22_X1 port map( A1 => n190, A2 => n64, B1 => n187, B2 => n126, ZN 
                           => n73);
   U37 : INV_X1 port map( A => i(4), ZN => n126);
   U38 : OAI22_X1 port map( A1 => n190, A2 => n63, B1 => n187, B2 => n125, ZN 
                           => n74);
   U39 : INV_X1 port map( A => i(5), ZN => n125);
   U40 : OAI22_X1 port map( A1 => n190, A2 => n62, B1 => n187, B2 => n124, ZN 
                           => n75);
   U41 : INV_X1 port map( A => i(6), ZN => n124);
   U42 : OAI22_X1 port map( A1 => n190, A2 => n61, B1 => n187, B2 => n123, ZN 
                           => n76);
   U43 : INV_X1 port map( A => i(7), ZN => n123);
   U44 : OAI22_X1 port map( A1 => n190, A2 => n60, B1 => n187, B2 => n122, ZN 
                           => n77);
   U45 : INV_X1 port map( A => i(8), ZN => n122);
   U46 : OAI22_X1 port map( A1 => n190, A2 => n59, B1 => n187, B2 => n121, ZN 
                           => n78);
   U47 : INV_X1 port map( A => i(9), ZN => n121);
   U48 : OAI22_X1 port map( A1 => n190, A2 => n58, B1 => n187, B2 => n120, ZN 
                           => n79);
   U49 : INV_X1 port map( A => i(10), ZN => n120);
   U50 : OAI22_X1 port map( A1 => n191, A2 => n57, B1 => n188, B2 => n119, ZN 
                           => n80);
   U51 : INV_X1 port map( A => i(11), ZN => n119);
   U52 : OAI22_X1 port map( A1 => n191, A2 => n56, B1 => n188, B2 => n118, ZN 
                           => n81);
   U53 : INV_X1 port map( A => i(12), ZN => n118);
   U54 : OAI22_X1 port map( A1 => n191, A2 => n55, B1 => n188, B2 => n117, ZN 
                           => n82);
   U55 : INV_X1 port map( A => i(13), ZN => n117);
   U56 : OAI22_X1 port map( A1 => n191, A2 => n54, B1 => n188, B2 => n116, ZN 
                           => n83);
   U57 : INV_X1 port map( A => i(14), ZN => n116);
   U58 : OAI22_X1 port map( A1 => n191, A2 => n53, B1 => n188, B2 => n115, ZN 
                           => n84);
   U59 : INV_X1 port map( A => i(15), ZN => n115);
   U60 : OAI22_X1 port map( A1 => n191, A2 => n52, B1 => n188, B2 => n114, ZN 
                           => n85);
   U61 : INV_X1 port map( A => i(16), ZN => n114);
   U62 : OAI22_X1 port map( A1 => n191, A2 => n51, B1 => n188, B2 => n113, ZN 
                           => n86);
   U63 : INV_X1 port map( A => i(17), ZN => n113);
   U64 : OAI22_X1 port map( A1 => n191, A2 => n50, B1 => n188, B2 => n112, ZN 
                           => n87);
   U65 : INV_X1 port map( A => i(18), ZN => n112);
   U66 : OAI22_X1 port map( A1 => n191, A2 => n49, B1 => n188, B2 => n111, ZN 
                           => n88);
   U67 : INV_X1 port map( A => i(19), ZN => n111);
   U68 : OAI22_X1 port map( A1 => n191, A2 => n48, B1 => n188, B2 => n110, ZN 
                           => n89);
   U69 : INV_X1 port map( A => i(20), ZN => n110);
   U70 : OAI22_X1 port map( A1 => n191, A2 => n47, B1 => n188, B2 => n109, ZN 
                           => n90);
   U71 : INV_X1 port map( A => i(21), ZN => n109);
   U72 : OAI22_X1 port map( A1 => n191, A2 => n46, B1 => n188, B2 => n108, ZN 
                           => n91);
   U73 : INV_X1 port map( A => i(22), ZN => n108);
   U74 : OAI22_X1 port map( A1 => n190, A2 => n37, B1 => n187, B2 => n131, ZN 
                           => n100);
   U75 : INV_X1 port map( A => i(31), ZN => n131);
   U76 : NAND2_X1 port map( A1 => n193, A2 => n190, ZN => n35);
   U77 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n34);
   U78 : INV_X1 port map( A => reset, ZN => n193);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity extensionModule26bit is

   port( i : in std_logic_vector (25 downto 0);  o : out std_logic_vector (31 
         downto 0));

end extensionModule26bit;

architecture SYN_Behavioral of extensionModule26bit is

begin
   o <= ( i(25), i(25), i(25), i(25), i(25), i(25), i(25), i(24), i(23), i(22),
      i(21), i(20), i(19), i(18), i(17), i(16), i(15), i(14), i(13), i(12), 
      i(11), i(10), i(9), i(8), i(7), i(6), i(5), i(4), i(3), i(2), i(1), i(0) 
      );

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity extensionModule is

   port( i : in std_logic_vector (15 downto 0);  o : out std_logic_vector (31 
         downto 0));

end extensionModule;

architecture SYN_Behavioral of extensionModule is

begin
   o <= ( i(15), i(15), i(15), i(15), i(15), i(15), i(15), i(15), i(15), i(15),
      i(15), i(15), i(15), i(15), i(15), i(15), i(15), i(14), i(13), i(12), 
      i(11), i(10), i(9), i(8), i(7), i(6), i(5), i(4), i(3), i(2), i(1), i(0) 
      );

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity register_file is

   port( data_in_port_w : in std_logic_vector (31 downto 0);  data_out_port_a, 
         data_out_port_b : out std_logic_vector (31 downto 0);  address_port_a,
         address_port_b, address_port_w : in std_logic_vector (4 downto 0);  
         r_signal_port_a, r_signal_port_b, w_signal, reset, enable : in 
         std_logic);

end register_file;

architecture SYN_Behavioral of register_file is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal registers_1_31_port, registers_1_30_port, registers_1_29_port, 
      registers_1_28_port, registers_1_27_port, registers_1_26_port, 
      registers_1_25_port, registers_1_24_port, registers_1_23_port, 
      registers_1_22_port, registers_1_21_port, registers_1_20_port, 
      registers_1_19_port, registers_1_18_port, registers_1_17_port, 
      registers_1_16_port, registers_1_15_port, registers_1_14_port, 
      registers_1_13_port, registers_1_12_port, registers_1_11_port, 
      registers_1_10_port, registers_1_9_port, registers_1_8_port, 
      registers_1_7_port, registers_1_6_port, registers_1_5_port, 
      registers_1_4_port, registers_1_3_port, registers_1_2_port, 
      registers_1_1_port, registers_1_0_port, registers_2_31_port, 
      registers_2_30_port, registers_2_29_port, registers_2_28_port, 
      registers_2_27_port, registers_2_26_port, registers_2_25_port, 
      registers_2_24_port, registers_2_23_port, registers_2_22_port, 
      registers_2_21_port, registers_2_20_port, registers_2_19_port, 
      registers_2_18_port, registers_2_17_port, registers_2_16_port, 
      registers_2_15_port, registers_2_14_port, registers_2_13_port, 
      registers_2_12_port, registers_2_11_port, registers_2_10_port, 
      registers_2_9_port, registers_2_8_port, registers_2_7_port, 
      registers_2_6_port, registers_2_5_port, registers_2_4_port, 
      registers_2_3_port, registers_2_2_port, registers_2_1_port, 
      registers_2_0_port, registers_3_31_port, registers_3_30_port, 
      registers_3_29_port, registers_3_28_port, registers_3_27_port, 
      registers_3_26_port, registers_3_25_port, registers_3_24_port, 
      registers_3_23_port, registers_3_22_port, registers_3_21_port, 
      registers_3_20_port, registers_3_19_port, registers_3_18_port, 
      registers_3_17_port, registers_3_16_port, registers_3_15_port, 
      registers_3_14_port, registers_3_13_port, registers_3_12_port, 
      registers_3_11_port, registers_3_10_port, registers_3_9_port, 
      registers_3_8_port, registers_3_7_port, registers_3_6_port, 
      registers_3_5_port, registers_3_4_port, registers_3_3_port, 
      registers_3_2_port, registers_3_1_port, registers_3_0_port, 
      registers_4_31_port, registers_4_30_port, registers_4_29_port, 
      registers_4_28_port, registers_4_27_port, registers_4_26_port, 
      registers_4_25_port, registers_4_24_port, registers_4_23_port, 
      registers_4_22_port, registers_4_21_port, registers_4_20_port, 
      registers_4_19_port, registers_4_18_port, registers_4_17_port, 
      registers_4_16_port, registers_4_15_port, registers_4_14_port, 
      registers_4_13_port, registers_4_12_port, registers_4_11_port, 
      registers_4_10_port, registers_4_9_port, registers_4_8_port, 
      registers_4_7_port, registers_4_6_port, registers_4_5_port, 
      registers_4_4_port, registers_4_3_port, registers_4_2_port, 
      registers_4_1_port, registers_4_0_port, registers_5_31_port, 
      registers_5_30_port, registers_5_29_port, registers_5_28_port, 
      registers_5_27_port, registers_5_26_port, registers_5_25_port, 
      registers_5_24_port, registers_5_23_port, registers_5_22_port, 
      registers_5_21_port, registers_5_20_port, registers_5_19_port, 
      registers_5_18_port, registers_5_17_port, registers_5_16_port, 
      registers_5_15_port, registers_5_14_port, registers_5_13_port, 
      registers_5_12_port, registers_5_11_port, registers_5_10_port, 
      registers_5_9_port, registers_5_8_port, registers_5_7_port, 
      registers_5_6_port, registers_5_5_port, registers_5_4_port, 
      registers_5_3_port, registers_5_2_port, registers_5_1_port, 
      registers_5_0_port, registers_6_31_port, registers_6_30_port, 
      registers_6_29_port, registers_6_28_port, registers_6_27_port, 
      registers_6_26_port, registers_6_25_port, registers_6_24_port, 
      registers_6_23_port, registers_6_22_port, registers_6_21_port, 
      registers_6_20_port, registers_6_19_port, registers_6_18_port, 
      registers_6_17_port, registers_6_16_port, registers_6_15_port, 
      registers_6_14_port, registers_6_13_port, registers_6_12_port, 
      registers_6_11_port, registers_6_10_port, registers_6_9_port, 
      registers_6_8_port, registers_6_7_port, registers_6_6_port, 
      registers_6_5_port, registers_6_4_port, registers_6_3_port, 
      registers_6_2_port, registers_6_1_port, registers_6_0_port, 
      registers_7_31_port, registers_7_30_port, registers_7_29_port, 
      registers_7_28_port, registers_7_27_port, registers_7_26_port, 
      registers_7_25_port, registers_7_24_port, registers_7_23_port, 
      registers_7_22_port, registers_7_21_port, registers_7_20_port, 
      registers_7_19_port, registers_7_18_port, registers_7_17_port, 
      registers_7_16_port, registers_7_15_port, registers_7_14_port, 
      registers_7_13_port, registers_7_12_port, registers_7_11_port, 
      registers_7_10_port, registers_7_9_port, registers_7_8_port, 
      registers_7_7_port, registers_7_6_port, registers_7_5_port, 
      registers_7_4_port, registers_7_3_port, registers_7_2_port, 
      registers_7_1_port, registers_7_0_port, registers_8_31_port, 
      registers_8_30_port, registers_8_29_port, registers_8_28_port, 
      registers_8_27_port, registers_8_26_port, registers_8_25_port, 
      registers_8_24_port, registers_8_23_port, registers_8_22_port, 
      registers_8_21_port, registers_8_20_port, registers_8_19_port, 
      registers_8_18_port, registers_8_17_port, registers_8_16_port, 
      registers_8_15_port, registers_8_14_port, registers_8_13_port, 
      registers_8_12_port, registers_8_11_port, registers_8_10_port, 
      registers_8_9_port, registers_8_8_port, registers_8_7_port, 
      registers_8_6_port, registers_8_5_port, registers_8_4_port, 
      registers_8_3_port, registers_8_2_port, registers_8_1_port, 
      registers_8_0_port, registers_9_31_port, registers_9_30_port, 
      registers_9_29_port, registers_9_28_port, registers_9_27_port, 
      registers_9_26_port, registers_9_25_port, registers_9_24_port, 
      registers_9_23_port, registers_9_22_port, registers_9_21_port, 
      registers_9_20_port, registers_9_19_port, registers_9_18_port, 
      registers_9_17_port, registers_9_16_port, registers_9_15_port, 
      registers_9_14_port, registers_9_13_port, registers_9_12_port, 
      registers_9_11_port, registers_9_10_port, registers_9_9_port, 
      registers_9_8_port, registers_9_7_port, registers_9_6_port, 
      registers_9_5_port, registers_9_4_port, registers_9_3_port, 
      registers_9_2_port, registers_9_1_port, registers_9_0_port, 
      registers_10_31_port, registers_10_30_port, registers_10_29_port, 
      registers_10_28_port, registers_10_27_port, registers_10_26_port, 
      registers_10_25_port, registers_10_24_port, registers_10_23_port, 
      registers_10_22_port, registers_10_21_port, registers_10_20_port, 
      registers_10_19_port, registers_10_18_port, registers_10_17_port, 
      registers_10_16_port, registers_10_15_port, registers_10_14_port, 
      registers_10_13_port, registers_10_12_port, registers_10_11_port, 
      registers_10_10_port, registers_10_9_port, registers_10_8_port, 
      registers_10_7_port, registers_10_6_port, registers_10_5_port, 
      registers_10_4_port, registers_10_3_port, registers_10_2_port, 
      registers_10_1_port, registers_10_0_port, registers_11_31_port, 
      registers_11_30_port, registers_11_29_port, registers_11_28_port, 
      registers_11_27_port, registers_11_26_port, registers_11_25_port, 
      registers_11_24_port, registers_11_23_port, registers_11_22_port, 
      registers_11_21_port, registers_11_20_port, registers_11_19_port, 
      registers_11_18_port, registers_11_17_port, registers_11_16_port, 
      registers_11_15_port, registers_11_14_port, registers_11_13_port, 
      registers_11_12_port, registers_11_11_port, registers_11_10_port, 
      registers_11_9_port, registers_11_8_port, registers_11_7_port, 
      registers_11_6_port, registers_11_5_port, registers_11_4_port, 
      registers_11_3_port, registers_11_2_port, registers_11_1_port, 
      registers_11_0_port, registers_12_31_port, registers_12_30_port, 
      registers_12_29_port, registers_12_28_port, registers_12_27_port, 
      registers_12_26_port, registers_12_25_port, registers_12_24_port, 
      registers_12_23_port, registers_12_22_port, registers_12_21_port, 
      registers_12_20_port, registers_12_19_port, registers_12_18_port, 
      registers_12_17_port, registers_12_16_port, registers_12_15_port, 
      registers_12_14_port, registers_12_13_port, registers_12_12_port, 
      registers_12_11_port, registers_12_10_port, registers_12_9_port, 
      registers_12_8_port, registers_12_7_port, registers_12_6_port, 
      registers_12_5_port, registers_12_4_port, registers_12_3_port, 
      registers_12_2_port, registers_12_1_port, registers_12_0_port, 
      registers_13_31_port, registers_13_30_port, registers_13_29_port, 
      registers_13_28_port, registers_13_27_port, registers_13_26_port, 
      registers_13_25_port, registers_13_24_port, registers_13_23_port, 
      registers_13_22_port, registers_13_21_port, registers_13_20_port, 
      registers_13_19_port, registers_13_18_port, registers_13_17_port, 
      registers_13_16_port, registers_13_15_port, registers_13_14_port, 
      registers_13_13_port, registers_13_12_port, registers_13_11_port, 
      registers_13_10_port, registers_13_9_port, registers_13_8_port, 
      registers_13_7_port, registers_13_6_port, registers_13_5_port, 
      registers_13_4_port, registers_13_3_port, registers_13_2_port, 
      registers_13_1_port, registers_13_0_port, registers_14_31_port, 
      registers_14_30_port, registers_14_29_port, registers_14_28_port, 
      registers_14_27_port, registers_14_26_port, registers_14_25_port, 
      registers_14_24_port, registers_14_23_port, registers_14_22_port, 
      registers_14_21_port, registers_14_20_port, registers_14_19_port, 
      registers_14_18_port, registers_14_17_port, registers_14_16_port, 
      registers_14_15_port, registers_14_14_port, registers_14_13_port, 
      registers_14_12_port, registers_14_11_port, registers_14_10_port, 
      registers_14_9_port, registers_14_8_port, registers_14_7_port, 
      registers_14_6_port, registers_14_5_port, registers_14_4_port, 
      registers_14_3_port, registers_14_2_port, registers_14_1_port, 
      registers_14_0_port, registers_15_31_port, registers_15_30_port, 
      registers_15_29_port, registers_15_28_port, registers_15_27_port, 
      registers_15_26_port, registers_15_25_port, registers_15_24_port, 
      registers_15_23_port, registers_15_22_port, registers_15_21_port, 
      registers_15_20_port, registers_15_19_port, registers_15_18_port, 
      registers_15_17_port, registers_15_16_port, registers_15_15_port, 
      registers_15_14_port, registers_15_13_port, registers_15_12_port, 
      registers_15_11_port, registers_15_10_port, registers_15_9_port, 
      registers_15_8_port, registers_15_7_port, registers_15_6_port, 
      registers_15_5_port, registers_15_4_port, registers_15_3_port, 
      registers_15_2_port, registers_15_1_port, registers_15_0_port, 
      registers_16_31_port, registers_16_30_port, registers_16_29_port, 
      registers_16_28_port, registers_16_27_port, registers_16_26_port, 
      registers_16_25_port, registers_16_24_port, registers_16_23_port, 
      registers_16_22_port, registers_16_21_port, registers_16_20_port, 
      registers_16_19_port, registers_16_18_port, registers_16_17_port, 
      registers_16_16_port, registers_16_15_port, registers_16_14_port, 
      registers_16_13_port, registers_16_12_port, registers_16_11_port, 
      registers_16_10_port, registers_16_9_port, registers_16_8_port, 
      registers_16_7_port, registers_16_6_port, registers_16_5_port, 
      registers_16_4_port, registers_16_3_port, registers_16_2_port, 
      registers_16_1_port, registers_16_0_port, registers_17_31_port, 
      registers_17_30_port, registers_17_29_port, registers_17_28_port, 
      registers_17_27_port, registers_17_26_port, registers_17_25_port, 
      registers_17_24_port, registers_17_23_port, registers_17_22_port, 
      registers_17_21_port, registers_17_20_port, registers_17_19_port, 
      registers_17_18_port, registers_17_17_port, registers_17_16_port, 
      registers_17_15_port, registers_17_14_port, registers_17_13_port, 
      registers_17_12_port, registers_17_11_port, registers_17_10_port, 
      registers_17_9_port, registers_17_8_port, registers_17_7_port, 
      registers_17_6_port, registers_17_5_port, registers_17_4_port, 
      registers_17_3_port, registers_17_2_port, registers_17_1_port, 
      registers_17_0_port, registers_18_31_port, registers_18_30_port, 
      registers_18_29_port, registers_18_28_port, registers_18_27_port, 
      registers_18_26_port, registers_18_25_port, registers_18_24_port, 
      registers_18_23_port, registers_18_22_port, registers_18_21_port, 
      registers_18_20_port, registers_18_19_port, registers_18_18_port, 
      registers_18_17_port, registers_18_16_port, registers_18_15_port, 
      registers_18_14_port, registers_18_13_port, registers_18_12_port, 
      registers_18_11_port, registers_18_10_port, registers_18_9_port, 
      registers_18_8_port, registers_18_7_port, registers_18_6_port, 
      registers_18_5_port, registers_18_4_port, registers_18_3_port, 
      registers_18_2_port, registers_18_1_port, registers_18_0_port, 
      registers_19_31_port, registers_19_30_port, registers_19_29_port, 
      registers_19_28_port, registers_19_27_port, registers_19_26_port, 
      registers_19_25_port, registers_19_24_port, registers_19_23_port, 
      registers_19_22_port, registers_19_21_port, registers_19_20_port, 
      registers_19_19_port, registers_19_18_port, registers_19_17_port, 
      registers_19_16_port, registers_19_15_port, registers_19_14_port, 
      registers_19_13_port, registers_19_12_port, registers_19_11_port, 
      registers_19_10_port, registers_19_9_port, registers_19_8_port, 
      registers_19_7_port, registers_19_6_port, registers_19_5_port, 
      registers_19_4_port, registers_19_3_port, registers_19_2_port, 
      registers_19_1_port, registers_19_0_port, registers_20_31_port, 
      registers_20_30_port, registers_20_29_port, registers_20_28_port, 
      registers_20_27_port, registers_20_26_port, registers_20_25_port, 
      registers_20_24_port, registers_20_23_port, registers_20_22_port, 
      registers_20_21_port, registers_20_20_port, registers_20_19_port, 
      registers_20_18_port, registers_20_17_port, registers_20_16_port, 
      registers_20_15_port, registers_20_14_port, registers_20_13_port, 
      registers_20_12_port, registers_20_11_port, registers_20_10_port, 
      registers_20_9_port, registers_20_8_port, registers_20_7_port, 
      registers_20_6_port, registers_20_5_port, registers_20_4_port, 
      registers_20_3_port, registers_20_2_port, registers_20_1_port, 
      registers_20_0_port, registers_21_31_port, registers_21_30_port, 
      registers_21_29_port, registers_21_28_port, registers_21_27_port, 
      registers_21_26_port, registers_21_25_port, registers_21_24_port, 
      registers_21_23_port, registers_21_22_port, registers_21_21_port, 
      registers_21_20_port, registers_21_19_port, registers_21_18_port, 
      registers_21_17_port, registers_21_16_port, registers_21_15_port, 
      registers_21_14_port, registers_21_13_port, registers_21_12_port, 
      registers_21_11_port, registers_21_10_port, registers_21_9_port, 
      registers_21_8_port, registers_21_7_port, registers_21_6_port, 
      registers_21_5_port, registers_21_4_port, registers_21_3_port, 
      registers_21_2_port, registers_21_1_port, registers_21_0_port, 
      registers_22_31_port, registers_22_30_port, registers_22_29_port, 
      registers_22_28_port, registers_22_27_port, registers_22_26_port, 
      registers_22_25_port, registers_22_24_port, registers_22_23_port, 
      registers_22_22_port, registers_22_21_port, registers_22_20_port, 
      registers_22_19_port, registers_22_18_port, registers_22_17_port, 
      registers_22_16_port, registers_22_15_port, registers_22_14_port, 
      registers_22_13_port, registers_22_12_port, registers_22_11_port, 
      registers_22_10_port, registers_22_9_port, registers_22_8_port, 
      registers_22_7_port, registers_22_6_port, registers_22_5_port, 
      registers_22_4_port, registers_22_3_port, registers_22_2_port, 
      registers_22_1_port, registers_22_0_port, registers_23_31_port, 
      registers_23_30_port, registers_23_29_port, registers_23_28_port, 
      registers_23_27_port, registers_23_26_port, registers_23_25_port, 
      registers_23_24_port, registers_23_23_port, registers_23_22_port, 
      registers_23_21_port, registers_23_20_port, registers_23_19_port, 
      registers_23_18_port, registers_23_17_port, registers_23_16_port, 
      registers_23_15_port, registers_23_14_port, registers_23_13_port, 
      registers_23_12_port, registers_23_11_port, registers_23_10_port, 
      registers_23_9_port, registers_23_8_port, registers_23_7_port, 
      registers_23_6_port, registers_23_5_port, registers_23_4_port, 
      registers_23_3_port, registers_23_2_port, registers_23_1_port, 
      registers_23_0_port, registers_24_31_port, registers_24_30_port, 
      registers_24_29_port, registers_24_28_port, registers_24_27_port, 
      registers_24_26_port, registers_24_25_port, registers_24_24_port, 
      registers_24_23_port, registers_24_22_port, registers_24_21_port, 
      registers_24_20_port, registers_24_19_port, registers_24_18_port, 
      registers_24_17_port, registers_24_16_port, registers_24_15_port, 
      registers_24_14_port, registers_24_13_port, registers_24_12_port, 
      registers_24_11_port, registers_24_10_port, registers_24_9_port, 
      registers_24_8_port, registers_24_7_port, registers_24_6_port, 
      registers_24_5_port, registers_24_4_port, registers_24_3_port, 
      registers_24_2_port, registers_24_1_port, registers_24_0_port, 
      registers_25_31_port, registers_25_30_port, registers_25_29_port, 
      registers_25_28_port, registers_25_27_port, registers_25_26_port, 
      registers_25_25_port, registers_25_24_port, registers_25_23_port, 
      registers_25_22_port, registers_25_21_port, registers_25_20_port, 
      registers_25_19_port, registers_25_18_port, registers_25_17_port, 
      registers_25_16_port, registers_25_15_port, registers_25_14_port, 
      registers_25_13_port, registers_25_12_port, registers_25_11_port, 
      registers_25_10_port, registers_25_9_port, registers_25_8_port, 
      registers_25_7_port, registers_25_6_port, registers_25_5_port, 
      registers_25_4_port, registers_25_3_port, registers_25_2_port, 
      registers_25_1_port, registers_25_0_port, registers_26_31_port, 
      registers_26_30_port, registers_26_29_port, registers_26_28_port, 
      registers_26_27_port, registers_26_26_port, registers_26_25_port, 
      registers_26_24_port, registers_26_23_port, registers_26_22_port, 
      registers_26_21_port, registers_26_20_port, registers_26_19_port, 
      registers_26_18_port, registers_26_17_port, registers_26_16_port, 
      registers_26_15_port, registers_26_14_port, registers_26_13_port, 
      registers_26_12_port, registers_26_11_port, registers_26_10_port, 
      registers_26_9_port, registers_26_8_port, registers_26_7_port, 
      registers_26_6_port, registers_26_5_port, registers_26_4_port, 
      registers_26_3_port, registers_26_2_port, registers_26_1_port, 
      registers_26_0_port, registers_27_31_port, registers_27_30_port, 
      registers_27_29_port, registers_27_28_port, registers_27_27_port, 
      registers_27_26_port, registers_27_25_port, registers_27_24_port, 
      registers_27_23_port, registers_27_22_port, registers_27_21_port, 
      registers_27_20_port, registers_27_19_port, registers_27_18_port, 
      registers_27_17_port, registers_27_16_port, registers_27_15_port, 
      registers_27_14_port, registers_27_13_port, registers_27_12_port, 
      registers_27_11_port, registers_27_10_port, registers_27_9_port, 
      registers_27_8_port, registers_27_7_port, registers_27_6_port, 
      registers_27_5_port, registers_27_4_port, registers_27_3_port, 
      registers_27_2_port, registers_27_1_port, registers_27_0_port, 
      registers_28_31_port, registers_28_30_port, registers_28_29_port, 
      registers_28_28_port, registers_28_27_port, registers_28_26_port, 
      registers_28_25_port, registers_28_24_port, registers_28_23_port, 
      registers_28_22_port, registers_28_21_port, registers_28_20_port, 
      registers_28_19_port, registers_28_18_port, registers_28_17_port, 
      registers_28_16_port, registers_28_15_port, registers_28_14_port, 
      registers_28_13_port, registers_28_12_port, registers_28_11_port, 
      registers_28_10_port, registers_28_9_port, registers_28_8_port, 
      registers_28_7_port, registers_28_6_port, registers_28_5_port, 
      registers_28_4_port, registers_28_3_port, registers_28_2_port, 
      registers_28_1_port, registers_28_0_port, registers_29_31_port, 
      registers_29_30_port, registers_29_29_port, registers_29_28_port, 
      registers_29_27_port, registers_29_26_port, registers_29_25_port, 
      registers_29_24_port, registers_29_23_port, registers_29_22_port, 
      registers_29_21_port, registers_29_20_port, registers_29_19_port, 
      registers_29_18_port, registers_29_17_port, registers_29_16_port, 
      registers_29_15_port, registers_29_14_port, registers_29_13_port, 
      registers_29_12_port, registers_29_11_port, registers_29_10_port, 
      registers_29_9_port, registers_29_8_port, registers_29_7_port, 
      registers_29_6_port, registers_29_5_port, registers_29_4_port, 
      registers_29_3_port, registers_29_2_port, registers_29_1_port, 
      registers_29_0_port, registers_30_31_port, registers_30_30_port, 
      registers_30_29_port, registers_30_28_port, registers_30_27_port, 
      registers_30_26_port, registers_30_25_port, registers_30_24_port, 
      registers_30_23_port, registers_30_22_port, registers_30_21_port, 
      registers_30_20_port, registers_30_19_port, registers_30_18_port, 
      registers_30_17_port, registers_30_16_port, registers_30_15_port, 
      registers_30_14_port, registers_30_13_port, registers_30_12_port, 
      registers_30_11_port, registers_30_10_port, registers_30_9_port, 
      registers_30_8_port, registers_30_7_port, registers_30_6_port, 
      registers_30_5_port, registers_30_4_port, registers_30_3_port, 
      registers_30_2_port, registers_30_1_port, registers_30_0_port, 
      registers_31_31_port, registers_31_30_port, registers_31_29_port, 
      registers_31_28_port, registers_31_27_port, registers_31_26_port, 
      registers_31_25_port, registers_31_24_port, registers_31_23_port, 
      registers_31_22_port, registers_31_21_port, registers_31_20_port, 
      registers_31_19_port, registers_31_18_port, registers_31_17_port, 
      registers_31_16_port, registers_31_15_port, registers_31_14_port, 
      registers_31_13_port, registers_31_12_port, registers_31_11_port, 
      registers_31_10_port, registers_31_9_port, registers_31_8_port, 
      registers_31_7_port, registers_31_6_port, registers_31_5_port, 
      registers_31_4_port, registers_31_3_port, registers_31_2_port, 
      registers_31_1_port, registers_31_0_port, n1778, n1779, n1780, n1781, 
      n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, 
      n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n2883, n2886, n2889, n2892, n2895, n2898, n2901, n2904, n2907, n2910, 
      n2913, n2916, n2919, n2922, n2925, n2928, n2931, n2934, n2937, n2940, 
      n2943, n2946, n2949, n2952, n2955, n2958, n2961, n2964, n2967, n2970, 
      n2973, n2976, n2979, n2982, n2985, n2988, n2991, n2994, n2997, n3000, 
      n3003, n3006, n3009, n3012, n3015, n3018, n3021, n3024, n3027, n3030, 
      n3033, n3036, n3039, n3042, n3045, n3048, n3051, n3054, n3057, n3060, 
      n3063, n3066, n3069, n3072, n3075, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1801, n1834, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, 
      n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, 
      n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, 
      n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, 
      n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, 
      n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, 
      n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, 
      n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, 
      n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, 
      n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, 
      n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, 
      n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, 
      n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, 
      n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, 
      n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, 
      n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, 
      n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, 
      n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, 
      n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, 
      n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, 
      n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, 
      n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, 
      n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, 
      n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, 
      n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, 
      n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, 
      n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, 
      n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, 
      n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, 
      n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, 
      n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, 
      n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, 
      n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
      n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, 
      n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, 
      n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, 
      n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, 
      n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, 
      n5176, n5177, n5178, n5179, n5180, n5181, n5182 : std_logic;

begin
   
   registers_reg_1_31_inst : DLH_X1 port map( G => n5086, D => n4989, Q => 
                           registers_1_31_port);
   registers_reg_1_30_inst : DLH_X1 port map( G => n5086, D => n4992, Q => 
                           registers_1_30_port);
   registers_reg_1_29_inst : DLH_X1 port map( G => n5086, D => n4995, Q => 
                           registers_1_29_port);
   registers_reg_1_28_inst : DLH_X1 port map( G => n5086, D => n4998, Q => 
                           registers_1_28_port);
   registers_reg_1_27_inst : DLH_X1 port map( G => n5086, D => n5001, Q => 
                           registers_1_27_port);
   registers_reg_1_26_inst : DLH_X1 port map( G => n5086, D => n5004, Q => 
                           registers_1_26_port);
   registers_reg_1_25_inst : DLH_X1 port map( G => n5086, D => n5007, Q => 
                           registers_1_25_port);
   registers_reg_1_24_inst : DLH_X1 port map( G => n5086, D => n5010, Q => 
                           registers_1_24_port);
   registers_reg_1_23_inst : DLH_X1 port map( G => n5086, D => n5013, Q => 
                           registers_1_23_port);
   registers_reg_1_22_inst : DLH_X1 port map( G => n5086, D => n5016, Q => 
                           registers_1_22_port);
   registers_reg_1_21_inst : DLH_X1 port map( G => n5085, D => n5019, Q => 
                           registers_1_21_port);
   registers_reg_1_20_inst : DLH_X1 port map( G => n5085, D => n5022, Q => 
                           registers_1_20_port);
   registers_reg_1_19_inst : DLH_X1 port map( G => n5085, D => n5025, Q => 
                           registers_1_19_port);
   registers_reg_1_18_inst : DLH_X1 port map( G => n5085, D => n5028, Q => 
                           registers_1_18_port);
   registers_reg_1_17_inst : DLH_X1 port map( G => n5085, D => n5031, Q => 
                           registers_1_17_port);
   registers_reg_1_16_inst : DLH_X1 port map( G => n5085, D => n5034, Q => 
                           registers_1_16_port);
   registers_reg_1_15_inst : DLH_X1 port map( G => n5085, D => n5037, Q => 
                           registers_1_15_port);
   registers_reg_1_14_inst : DLH_X1 port map( G => n5085, D => n5040, Q => 
                           registers_1_14_port);
   registers_reg_1_13_inst : DLH_X1 port map( G => n5085, D => n5043, Q => 
                           registers_1_13_port);
   registers_reg_1_12_inst : DLH_X1 port map( G => n5085, D => n5046, Q => 
                           registers_1_12_port);
   registers_reg_1_11_inst : DLH_X1 port map( G => n5085, D => n5049, Q => 
                           registers_1_11_port);
   registers_reg_1_10_inst : DLH_X1 port map( G => n5084, D => n5052, Q => 
                           registers_1_10_port);
   registers_reg_1_9_inst : DLH_X1 port map( G => n5084, D => n5055, Q => 
                           registers_1_9_port);
   registers_reg_1_8_inst : DLH_X1 port map( G => n5084, D => n5058, Q => 
                           registers_1_8_port);
   registers_reg_1_7_inst : DLH_X1 port map( G => n5084, D => n5061, Q => 
                           registers_1_7_port);
   registers_reg_1_6_inst : DLH_X1 port map( G => n5084, D => n5064, Q => 
                           registers_1_6_port);
   registers_reg_1_5_inst : DLH_X1 port map( G => n5084, D => n5067, Q => 
                           registers_1_5_port);
   registers_reg_1_4_inst : DLH_X1 port map( G => n5084, D => n5070, Q => 
                           registers_1_4_port);
   registers_reg_1_3_inst : DLH_X1 port map( G => n5084, D => n5073, Q => 
                           registers_1_3_port);
   registers_reg_1_2_inst : DLH_X1 port map( G => n5084, D => n5076, Q => 
                           registers_1_2_port);
   registers_reg_1_1_inst : DLH_X1 port map( G => n5084, D => n5079, Q => 
                           registers_1_1_port);
   registers_reg_1_0_inst : DLH_X1 port map( G => n5084, D => n5082, Q => 
                           registers_1_0_port);
   registers_reg_2_31_inst : DLH_X1 port map( G => n5089, D => n4989, Q => 
                           registers_2_31_port);
   registers_reg_2_30_inst : DLH_X1 port map( G => n5089, D => n4992, Q => 
                           registers_2_30_port);
   registers_reg_2_29_inst : DLH_X1 port map( G => n5089, D => n4995, Q => 
                           registers_2_29_port);
   registers_reg_2_28_inst : DLH_X1 port map( G => n5089, D => n4998, Q => 
                           registers_2_28_port);
   registers_reg_2_27_inst : DLH_X1 port map( G => n5089, D => n5001, Q => 
                           registers_2_27_port);
   registers_reg_2_26_inst : DLH_X1 port map( G => n5089, D => n5004, Q => 
                           registers_2_26_port);
   registers_reg_2_25_inst : DLH_X1 port map( G => n5089, D => n5007, Q => 
                           registers_2_25_port);
   registers_reg_2_24_inst : DLH_X1 port map( G => n5089, D => n5010, Q => 
                           registers_2_24_port);
   registers_reg_2_23_inst : DLH_X1 port map( G => n5089, D => n5013, Q => 
                           registers_2_23_port);
   registers_reg_2_22_inst : DLH_X1 port map( G => n5089, D => n5016, Q => 
                           registers_2_22_port);
   registers_reg_2_21_inst : DLH_X1 port map( G => n5088, D => n5019, Q => 
                           registers_2_21_port);
   registers_reg_2_20_inst : DLH_X1 port map( G => n5088, D => n5022, Q => 
                           registers_2_20_port);
   registers_reg_2_19_inst : DLH_X1 port map( G => n5088, D => n5025, Q => 
                           registers_2_19_port);
   registers_reg_2_18_inst : DLH_X1 port map( G => n5088, D => n5028, Q => 
                           registers_2_18_port);
   registers_reg_2_17_inst : DLH_X1 port map( G => n5088, D => n5031, Q => 
                           registers_2_17_port);
   registers_reg_2_16_inst : DLH_X1 port map( G => n5088, D => n5034, Q => 
                           registers_2_16_port);
   registers_reg_2_15_inst : DLH_X1 port map( G => n5088, D => n5037, Q => 
                           registers_2_15_port);
   registers_reg_2_14_inst : DLH_X1 port map( G => n5088, D => n5040, Q => 
                           registers_2_14_port);
   registers_reg_2_13_inst : DLH_X1 port map( G => n5088, D => n5043, Q => 
                           registers_2_13_port);
   registers_reg_2_12_inst : DLH_X1 port map( G => n5088, D => n5046, Q => 
                           registers_2_12_port);
   registers_reg_2_11_inst : DLH_X1 port map( G => n5088, D => n5049, Q => 
                           registers_2_11_port);
   registers_reg_2_10_inst : DLH_X1 port map( G => n5087, D => n5052, Q => 
                           registers_2_10_port);
   registers_reg_2_9_inst : DLH_X1 port map( G => n5087, D => n5055, Q => 
                           registers_2_9_port);
   registers_reg_2_8_inst : DLH_X1 port map( G => n5087, D => n5058, Q => 
                           registers_2_8_port);
   registers_reg_2_7_inst : DLH_X1 port map( G => n5087, D => n5061, Q => 
                           registers_2_7_port);
   registers_reg_2_6_inst : DLH_X1 port map( G => n5087, D => n5064, Q => 
                           registers_2_6_port);
   registers_reg_2_5_inst : DLH_X1 port map( G => n5087, D => n5067, Q => 
                           registers_2_5_port);
   registers_reg_2_4_inst : DLH_X1 port map( G => n5087, D => n5070, Q => 
                           registers_2_4_port);
   registers_reg_2_3_inst : DLH_X1 port map( G => n5087, D => n5073, Q => 
                           registers_2_3_port);
   registers_reg_2_2_inst : DLH_X1 port map( G => n5087, D => n5076, Q => 
                           registers_2_2_port);
   registers_reg_2_1_inst : DLH_X1 port map( G => n5087, D => n5079, Q => 
                           registers_2_1_port);
   registers_reg_2_0_inst : DLH_X1 port map( G => n5087, D => n5082, Q => 
                           registers_2_0_port);
   registers_reg_3_31_inst : DLH_X1 port map( G => n5092, D => n4990, Q => 
                           registers_3_31_port);
   registers_reg_3_30_inst : DLH_X1 port map( G => n5092, D => n4993, Q => 
                           registers_3_30_port);
   registers_reg_3_29_inst : DLH_X1 port map( G => n5092, D => n4996, Q => 
                           registers_3_29_port);
   registers_reg_3_28_inst : DLH_X1 port map( G => n5092, D => n4999, Q => 
                           registers_3_28_port);
   registers_reg_3_27_inst : DLH_X1 port map( G => n5092, D => n5002, Q => 
                           registers_3_27_port);
   registers_reg_3_26_inst : DLH_X1 port map( G => n5092, D => n5005, Q => 
                           registers_3_26_port);
   registers_reg_3_25_inst : DLH_X1 port map( G => n5092, D => n5008, Q => 
                           registers_3_25_port);
   registers_reg_3_24_inst : DLH_X1 port map( G => n5092, D => n5011, Q => 
                           registers_3_24_port);
   registers_reg_3_23_inst : DLH_X1 port map( G => n5092, D => n5014, Q => 
                           registers_3_23_port);
   registers_reg_3_22_inst : DLH_X1 port map( G => n5092, D => n5017, Q => 
                           registers_3_22_port);
   registers_reg_3_21_inst : DLH_X1 port map( G => n5091, D => n5020, Q => 
                           registers_3_21_port);
   registers_reg_3_20_inst : DLH_X1 port map( G => n5091, D => n5023, Q => 
                           registers_3_20_port);
   registers_reg_3_19_inst : DLH_X1 port map( G => n5091, D => n5026, Q => 
                           registers_3_19_port);
   registers_reg_3_18_inst : DLH_X1 port map( G => n5091, D => n5029, Q => 
                           registers_3_18_port);
   registers_reg_3_17_inst : DLH_X1 port map( G => n5091, D => n5032, Q => 
                           registers_3_17_port);
   registers_reg_3_16_inst : DLH_X1 port map( G => n5091, D => n5035, Q => 
                           registers_3_16_port);
   registers_reg_3_15_inst : DLH_X1 port map( G => n5091, D => n5038, Q => 
                           registers_3_15_port);
   registers_reg_3_14_inst : DLH_X1 port map( G => n5091, D => n5041, Q => 
                           registers_3_14_port);
   registers_reg_3_13_inst : DLH_X1 port map( G => n5091, D => n5044, Q => 
                           registers_3_13_port);
   registers_reg_3_12_inst : DLH_X1 port map( G => n5091, D => n5047, Q => 
                           registers_3_12_port);
   registers_reg_3_11_inst : DLH_X1 port map( G => n5091, D => n5050, Q => 
                           registers_3_11_port);
   registers_reg_3_10_inst : DLH_X1 port map( G => n5090, D => n5053, Q => 
                           registers_3_10_port);
   registers_reg_3_9_inst : DLH_X1 port map( G => n5090, D => n5056, Q => 
                           registers_3_9_port);
   registers_reg_3_8_inst : DLH_X1 port map( G => n5090, D => n5059, Q => 
                           registers_3_8_port);
   registers_reg_3_7_inst : DLH_X1 port map( G => n5090, D => n5062, Q => 
                           registers_3_7_port);
   registers_reg_3_6_inst : DLH_X1 port map( G => n5090, D => n5065, Q => 
                           registers_3_6_port);
   registers_reg_3_5_inst : DLH_X1 port map( G => n5090, D => n5068, Q => 
                           registers_3_5_port);
   registers_reg_3_4_inst : DLH_X1 port map( G => n5090, D => n5071, Q => 
                           registers_3_4_port);
   registers_reg_3_3_inst : DLH_X1 port map( G => n5090, D => n5074, Q => 
                           registers_3_3_port);
   registers_reg_3_2_inst : DLH_X1 port map( G => n5090, D => n5077, Q => 
                           registers_3_2_port);
   registers_reg_3_1_inst : DLH_X1 port map( G => n5090, D => n5080, Q => 
                           registers_3_1_port);
   registers_reg_3_0_inst : DLH_X1 port map( G => n5090, D => n5083, Q => 
                           registers_3_0_port);
   registers_reg_4_31_inst : DLH_X1 port map( G => n5095, D => n4990, Q => 
                           registers_4_31_port);
   registers_reg_4_30_inst : DLH_X1 port map( G => n5095, D => n4993, Q => 
                           registers_4_30_port);
   registers_reg_4_29_inst : DLH_X1 port map( G => n5095, D => n4996, Q => 
                           registers_4_29_port);
   registers_reg_4_28_inst : DLH_X1 port map( G => n5095, D => n4999, Q => 
                           registers_4_28_port);
   registers_reg_4_27_inst : DLH_X1 port map( G => n5095, D => n5002, Q => 
                           registers_4_27_port);
   registers_reg_4_26_inst : DLH_X1 port map( G => n5095, D => n5005, Q => 
                           registers_4_26_port);
   registers_reg_4_25_inst : DLH_X1 port map( G => n5095, D => n5008, Q => 
                           registers_4_25_port);
   registers_reg_4_24_inst : DLH_X1 port map( G => n5095, D => n5011, Q => 
                           registers_4_24_port);
   registers_reg_4_23_inst : DLH_X1 port map( G => n5095, D => n5014, Q => 
                           registers_4_23_port);
   registers_reg_4_22_inst : DLH_X1 port map( G => n5095, D => n5017, Q => 
                           registers_4_22_port);
   registers_reg_4_21_inst : DLH_X1 port map( G => n5094, D => n5020, Q => 
                           registers_4_21_port);
   registers_reg_4_20_inst : DLH_X1 port map( G => n5094, D => n5023, Q => 
                           registers_4_20_port);
   registers_reg_4_19_inst : DLH_X1 port map( G => n5094, D => n5026, Q => 
                           registers_4_19_port);
   registers_reg_4_18_inst : DLH_X1 port map( G => n5094, D => n5029, Q => 
                           registers_4_18_port);
   registers_reg_4_17_inst : DLH_X1 port map( G => n5094, D => n5032, Q => 
                           registers_4_17_port);
   registers_reg_4_16_inst : DLH_X1 port map( G => n5094, D => n5035, Q => 
                           registers_4_16_port);
   registers_reg_4_15_inst : DLH_X1 port map( G => n5094, D => n5038, Q => 
                           registers_4_15_port);
   registers_reg_4_14_inst : DLH_X1 port map( G => n5094, D => n5041, Q => 
                           registers_4_14_port);
   registers_reg_4_13_inst : DLH_X1 port map( G => n5094, D => n5044, Q => 
                           registers_4_13_port);
   registers_reg_4_12_inst : DLH_X1 port map( G => n5094, D => n5047, Q => 
                           registers_4_12_port);
   registers_reg_4_11_inst : DLH_X1 port map( G => n5094, D => n5050, Q => 
                           registers_4_11_port);
   registers_reg_4_10_inst : DLH_X1 port map( G => n5093, D => n5053, Q => 
                           registers_4_10_port);
   registers_reg_4_9_inst : DLH_X1 port map( G => n5093, D => n5056, Q => 
                           registers_4_9_port);
   registers_reg_4_8_inst : DLH_X1 port map( G => n5093, D => n5059, Q => 
                           registers_4_8_port);
   registers_reg_4_7_inst : DLH_X1 port map( G => n5093, D => n5062, Q => 
                           registers_4_7_port);
   registers_reg_4_6_inst : DLH_X1 port map( G => n5093, D => n5065, Q => 
                           registers_4_6_port);
   registers_reg_4_5_inst : DLH_X1 port map( G => n5093, D => n5068, Q => 
                           registers_4_5_port);
   registers_reg_4_4_inst : DLH_X1 port map( G => n5093, D => n5071, Q => 
                           registers_4_4_port);
   registers_reg_4_3_inst : DLH_X1 port map( G => n5093, D => n5074, Q => 
                           registers_4_3_port);
   registers_reg_4_2_inst : DLH_X1 port map( G => n5093, D => n5077, Q => 
                           registers_4_2_port);
   registers_reg_4_1_inst : DLH_X1 port map( G => n5093, D => n5080, Q => 
                           registers_4_1_port);
   registers_reg_4_0_inst : DLH_X1 port map( G => n5093, D => n5083, Q => 
                           registers_4_0_port);
   registers_reg_5_31_inst : DLH_X1 port map( G => n5098, D => n4990, Q => 
                           registers_5_31_port);
   registers_reg_5_30_inst : DLH_X1 port map( G => n5098, D => n4993, Q => 
                           registers_5_30_port);
   registers_reg_5_29_inst : DLH_X1 port map( G => n5098, D => n4996, Q => 
                           registers_5_29_port);
   registers_reg_5_28_inst : DLH_X1 port map( G => n5098, D => n4999, Q => 
                           registers_5_28_port);
   registers_reg_5_27_inst : DLH_X1 port map( G => n5098, D => n5002, Q => 
                           registers_5_27_port);
   registers_reg_5_26_inst : DLH_X1 port map( G => n5098, D => n5005, Q => 
                           registers_5_26_port);
   registers_reg_5_25_inst : DLH_X1 port map( G => n5098, D => n5008, Q => 
                           registers_5_25_port);
   registers_reg_5_24_inst : DLH_X1 port map( G => n5098, D => n5011, Q => 
                           registers_5_24_port);
   registers_reg_5_23_inst : DLH_X1 port map( G => n5098, D => n5014, Q => 
                           registers_5_23_port);
   registers_reg_5_22_inst : DLH_X1 port map( G => n5098, D => n5017, Q => 
                           registers_5_22_port);
   registers_reg_5_21_inst : DLH_X1 port map( G => n5097, D => n5020, Q => 
                           registers_5_21_port);
   registers_reg_5_20_inst : DLH_X1 port map( G => n5097, D => n5023, Q => 
                           registers_5_20_port);
   registers_reg_5_19_inst : DLH_X1 port map( G => n5097, D => n5026, Q => 
                           registers_5_19_port);
   registers_reg_5_18_inst : DLH_X1 port map( G => n5097, D => n5029, Q => 
                           registers_5_18_port);
   registers_reg_5_17_inst : DLH_X1 port map( G => n5097, D => n5032, Q => 
                           registers_5_17_port);
   registers_reg_5_16_inst : DLH_X1 port map( G => n5097, D => n5035, Q => 
                           registers_5_16_port);
   registers_reg_5_15_inst : DLH_X1 port map( G => n5097, D => n5038, Q => 
                           registers_5_15_port);
   registers_reg_5_14_inst : DLH_X1 port map( G => n5097, D => n5041, Q => 
                           registers_5_14_port);
   registers_reg_5_13_inst : DLH_X1 port map( G => n5097, D => n5044, Q => 
                           registers_5_13_port);
   registers_reg_5_12_inst : DLH_X1 port map( G => n5097, D => n5047, Q => 
                           registers_5_12_port);
   registers_reg_5_11_inst : DLH_X1 port map( G => n5097, D => n5050, Q => 
                           registers_5_11_port);
   registers_reg_5_10_inst : DLH_X1 port map( G => n5096, D => n5053, Q => 
                           registers_5_10_port);
   registers_reg_5_9_inst : DLH_X1 port map( G => n5096, D => n5056, Q => 
                           registers_5_9_port);
   registers_reg_5_8_inst : DLH_X1 port map( G => n5096, D => n5059, Q => 
                           registers_5_8_port);
   registers_reg_5_7_inst : DLH_X1 port map( G => n5096, D => n5062, Q => 
                           registers_5_7_port);
   registers_reg_5_6_inst : DLH_X1 port map( G => n5096, D => n5065, Q => 
                           registers_5_6_port);
   registers_reg_5_5_inst : DLH_X1 port map( G => n5096, D => n5068, Q => 
                           registers_5_5_port);
   registers_reg_5_4_inst : DLH_X1 port map( G => n5096, D => n5071, Q => 
                           registers_5_4_port);
   registers_reg_5_3_inst : DLH_X1 port map( G => n5096, D => n5074, Q => 
                           registers_5_3_port);
   registers_reg_5_2_inst : DLH_X1 port map( G => n5096, D => n5077, Q => 
                           registers_5_2_port);
   registers_reg_5_1_inst : DLH_X1 port map( G => n5096, D => n5080, Q => 
                           registers_5_1_port);
   registers_reg_5_0_inst : DLH_X1 port map( G => n5096, D => n5083, Q => 
                           registers_5_0_port);
   registers_reg_6_31_inst : DLH_X1 port map( G => n5101, D => n4990, Q => 
                           registers_6_31_port);
   registers_reg_6_30_inst : DLH_X1 port map( G => n5101, D => n4993, Q => 
                           registers_6_30_port);
   registers_reg_6_29_inst : DLH_X1 port map( G => n5101, D => n4996, Q => 
                           registers_6_29_port);
   registers_reg_6_28_inst : DLH_X1 port map( G => n5101, D => n4999, Q => 
                           registers_6_28_port);
   registers_reg_6_27_inst : DLH_X1 port map( G => n5101, D => n5002, Q => 
                           registers_6_27_port);
   registers_reg_6_26_inst : DLH_X1 port map( G => n5101, D => n5005, Q => 
                           registers_6_26_port);
   registers_reg_6_25_inst : DLH_X1 port map( G => n5101, D => n5008, Q => 
                           registers_6_25_port);
   registers_reg_6_24_inst : DLH_X1 port map( G => n5101, D => n5011, Q => 
                           registers_6_24_port);
   registers_reg_6_23_inst : DLH_X1 port map( G => n5101, D => n5014, Q => 
                           registers_6_23_port);
   registers_reg_6_22_inst : DLH_X1 port map( G => n5101, D => n5017, Q => 
                           registers_6_22_port);
   registers_reg_6_21_inst : DLH_X1 port map( G => n5100, D => n5020, Q => 
                           registers_6_21_port);
   registers_reg_6_20_inst : DLH_X1 port map( G => n5100, D => n5023, Q => 
                           registers_6_20_port);
   registers_reg_6_19_inst : DLH_X1 port map( G => n5100, D => n5026, Q => 
                           registers_6_19_port);
   registers_reg_6_18_inst : DLH_X1 port map( G => n5100, D => n5029, Q => 
                           registers_6_18_port);
   registers_reg_6_17_inst : DLH_X1 port map( G => n5100, D => n5032, Q => 
                           registers_6_17_port);
   registers_reg_6_16_inst : DLH_X1 port map( G => n5100, D => n5035, Q => 
                           registers_6_16_port);
   registers_reg_6_15_inst : DLH_X1 port map( G => n5100, D => n5038, Q => 
                           registers_6_15_port);
   registers_reg_6_14_inst : DLH_X1 port map( G => n5100, D => n5041, Q => 
                           registers_6_14_port);
   registers_reg_6_13_inst : DLH_X1 port map( G => n5100, D => n5044, Q => 
                           registers_6_13_port);
   registers_reg_6_12_inst : DLH_X1 port map( G => n5100, D => n5047, Q => 
                           registers_6_12_port);
   registers_reg_6_11_inst : DLH_X1 port map( G => n5100, D => n5050, Q => 
                           registers_6_11_port);
   registers_reg_6_10_inst : DLH_X1 port map( G => n5099, D => n5053, Q => 
                           registers_6_10_port);
   registers_reg_6_9_inst : DLH_X1 port map( G => n5099, D => n5056, Q => 
                           registers_6_9_port);
   registers_reg_6_8_inst : DLH_X1 port map( G => n5099, D => n5059, Q => 
                           registers_6_8_port);
   registers_reg_6_7_inst : DLH_X1 port map( G => n5099, D => n5062, Q => 
                           registers_6_7_port);
   registers_reg_6_6_inst : DLH_X1 port map( G => n5099, D => n5065, Q => 
                           registers_6_6_port);
   registers_reg_6_5_inst : DLH_X1 port map( G => n5099, D => n5068, Q => 
                           registers_6_5_port);
   registers_reg_6_4_inst : DLH_X1 port map( G => n5099, D => n5071, Q => 
                           registers_6_4_port);
   registers_reg_6_3_inst : DLH_X1 port map( G => n5099, D => n5074, Q => 
                           registers_6_3_port);
   registers_reg_6_2_inst : DLH_X1 port map( G => n5099, D => n5077, Q => 
                           registers_6_2_port);
   registers_reg_6_1_inst : DLH_X1 port map( G => n5099, D => n5080, Q => 
                           registers_6_1_port);
   registers_reg_6_0_inst : DLH_X1 port map( G => n5099, D => n5083, Q => 
                           registers_6_0_port);
   registers_reg_7_31_inst : DLH_X1 port map( G => n5104, D => n4990, Q => 
                           registers_7_31_port);
   registers_reg_7_30_inst : DLH_X1 port map( G => n5104, D => n4993, Q => 
                           registers_7_30_port);
   registers_reg_7_29_inst : DLH_X1 port map( G => n5104, D => n4996, Q => 
                           registers_7_29_port);
   registers_reg_7_28_inst : DLH_X1 port map( G => n5104, D => n4999, Q => 
                           registers_7_28_port);
   registers_reg_7_27_inst : DLH_X1 port map( G => n5104, D => n5002, Q => 
                           registers_7_27_port);
   registers_reg_7_26_inst : DLH_X1 port map( G => n5104, D => n5005, Q => 
                           registers_7_26_port);
   registers_reg_7_25_inst : DLH_X1 port map( G => n5104, D => n5008, Q => 
                           registers_7_25_port);
   registers_reg_7_24_inst : DLH_X1 port map( G => n5104, D => n5011, Q => 
                           registers_7_24_port);
   registers_reg_7_23_inst : DLH_X1 port map( G => n5104, D => n5014, Q => 
                           registers_7_23_port);
   registers_reg_7_22_inst : DLH_X1 port map( G => n5104, D => n5017, Q => 
                           registers_7_22_port);
   registers_reg_7_21_inst : DLH_X1 port map( G => n5103, D => n5020, Q => 
                           registers_7_21_port);
   registers_reg_7_20_inst : DLH_X1 port map( G => n5103, D => n5023, Q => 
                           registers_7_20_port);
   registers_reg_7_19_inst : DLH_X1 port map( G => n5103, D => n5026, Q => 
                           registers_7_19_port);
   registers_reg_7_18_inst : DLH_X1 port map( G => n5103, D => n5029, Q => 
                           registers_7_18_port);
   registers_reg_7_17_inst : DLH_X1 port map( G => n5103, D => n5032, Q => 
                           registers_7_17_port);
   registers_reg_7_16_inst : DLH_X1 port map( G => n5103, D => n5035, Q => 
                           registers_7_16_port);
   registers_reg_7_15_inst : DLH_X1 port map( G => n5103, D => n5038, Q => 
                           registers_7_15_port);
   registers_reg_7_14_inst : DLH_X1 port map( G => n5103, D => n5041, Q => 
                           registers_7_14_port);
   registers_reg_7_13_inst : DLH_X1 port map( G => n5103, D => n5044, Q => 
                           registers_7_13_port);
   registers_reg_7_12_inst : DLH_X1 port map( G => n5103, D => n5047, Q => 
                           registers_7_12_port);
   registers_reg_7_11_inst : DLH_X1 port map( G => n5103, D => n5050, Q => 
                           registers_7_11_port);
   registers_reg_7_10_inst : DLH_X1 port map( G => n5102, D => n5053, Q => 
                           registers_7_10_port);
   registers_reg_7_9_inst : DLH_X1 port map( G => n5102, D => n5056, Q => 
                           registers_7_9_port);
   registers_reg_7_8_inst : DLH_X1 port map( G => n5102, D => n5059, Q => 
                           registers_7_8_port);
   registers_reg_7_7_inst : DLH_X1 port map( G => n5102, D => n5062, Q => 
                           registers_7_7_port);
   registers_reg_7_6_inst : DLH_X1 port map( G => n5102, D => n5065, Q => 
                           registers_7_6_port);
   registers_reg_7_5_inst : DLH_X1 port map( G => n5102, D => n5068, Q => 
                           registers_7_5_port);
   registers_reg_7_4_inst : DLH_X1 port map( G => n5102, D => n5071, Q => 
                           registers_7_4_port);
   registers_reg_7_3_inst : DLH_X1 port map( G => n5102, D => n5074, Q => 
                           registers_7_3_port);
   registers_reg_7_2_inst : DLH_X1 port map( G => n5102, D => n5077, Q => 
                           registers_7_2_port);
   registers_reg_7_1_inst : DLH_X1 port map( G => n5102, D => n5080, Q => 
                           registers_7_1_port);
   registers_reg_7_0_inst : DLH_X1 port map( G => n5102, D => n5083, Q => 
                           registers_7_0_port);
   registers_reg_8_31_inst : DLH_X1 port map( G => n5107, D => n4990, Q => 
                           registers_8_31_port);
   registers_reg_8_30_inst : DLH_X1 port map( G => n5107, D => n4993, Q => 
                           registers_8_30_port);
   registers_reg_8_29_inst : DLH_X1 port map( G => n5107, D => n4996, Q => 
                           registers_8_29_port);
   registers_reg_8_28_inst : DLH_X1 port map( G => n5107, D => n4999, Q => 
                           registers_8_28_port);
   registers_reg_8_27_inst : DLH_X1 port map( G => n5107, D => n5002, Q => 
                           registers_8_27_port);
   registers_reg_8_26_inst : DLH_X1 port map( G => n5107, D => n5005, Q => 
                           registers_8_26_port);
   registers_reg_8_25_inst : DLH_X1 port map( G => n5107, D => n5008, Q => 
                           registers_8_25_port);
   registers_reg_8_24_inst : DLH_X1 port map( G => n5107, D => n5011, Q => 
                           registers_8_24_port);
   registers_reg_8_23_inst : DLH_X1 port map( G => n5107, D => n5014, Q => 
                           registers_8_23_port);
   registers_reg_8_22_inst : DLH_X1 port map( G => n5107, D => n5017, Q => 
                           registers_8_22_port);
   registers_reg_8_21_inst : DLH_X1 port map( G => n5106, D => n5020, Q => 
                           registers_8_21_port);
   registers_reg_8_20_inst : DLH_X1 port map( G => n5106, D => n5023, Q => 
                           registers_8_20_port);
   registers_reg_8_19_inst : DLH_X1 port map( G => n5106, D => n5026, Q => 
                           registers_8_19_port);
   registers_reg_8_18_inst : DLH_X1 port map( G => n5106, D => n5029, Q => 
                           registers_8_18_port);
   registers_reg_8_17_inst : DLH_X1 port map( G => n5106, D => n5032, Q => 
                           registers_8_17_port);
   registers_reg_8_16_inst : DLH_X1 port map( G => n5106, D => n5035, Q => 
                           registers_8_16_port);
   registers_reg_8_15_inst : DLH_X1 port map( G => n5106, D => n5038, Q => 
                           registers_8_15_port);
   registers_reg_8_14_inst : DLH_X1 port map( G => n5106, D => n5041, Q => 
                           registers_8_14_port);
   registers_reg_8_13_inst : DLH_X1 port map( G => n5106, D => n5044, Q => 
                           registers_8_13_port);
   registers_reg_8_12_inst : DLH_X1 port map( G => n5106, D => n5047, Q => 
                           registers_8_12_port);
   registers_reg_8_11_inst : DLH_X1 port map( G => n5106, D => n5050, Q => 
                           registers_8_11_port);
   registers_reg_8_10_inst : DLH_X1 port map( G => n5105, D => n5053, Q => 
                           registers_8_10_port);
   registers_reg_8_9_inst : DLH_X1 port map( G => n5105, D => n5056, Q => 
                           registers_8_9_port);
   registers_reg_8_8_inst : DLH_X1 port map( G => n5105, D => n5059, Q => 
                           registers_8_8_port);
   registers_reg_8_7_inst : DLH_X1 port map( G => n5105, D => n5062, Q => 
                           registers_8_7_port);
   registers_reg_8_6_inst : DLH_X1 port map( G => n5105, D => n5065, Q => 
                           registers_8_6_port);
   registers_reg_8_5_inst : DLH_X1 port map( G => n5105, D => n5068, Q => 
                           registers_8_5_port);
   registers_reg_8_4_inst : DLH_X1 port map( G => n5105, D => n5071, Q => 
                           registers_8_4_port);
   registers_reg_8_3_inst : DLH_X1 port map( G => n5105, D => n5074, Q => 
                           registers_8_3_port);
   registers_reg_8_2_inst : DLH_X1 port map( G => n5105, D => n5077, Q => 
                           registers_8_2_port);
   registers_reg_8_1_inst : DLH_X1 port map( G => n5105, D => n5080, Q => 
                           registers_8_1_port);
   registers_reg_8_0_inst : DLH_X1 port map( G => n5105, D => n5083, Q => 
                           registers_8_0_port);
   registers_reg_9_31_inst : DLH_X1 port map( G => n5110, D => n4990, Q => 
                           registers_9_31_port);
   registers_reg_9_30_inst : DLH_X1 port map( G => n5110, D => n4993, Q => 
                           registers_9_30_port);
   registers_reg_9_29_inst : DLH_X1 port map( G => n5110, D => n4996, Q => 
                           registers_9_29_port);
   registers_reg_9_28_inst : DLH_X1 port map( G => n5110, D => n4999, Q => 
                           registers_9_28_port);
   registers_reg_9_27_inst : DLH_X1 port map( G => n5110, D => n5002, Q => 
                           registers_9_27_port);
   registers_reg_9_26_inst : DLH_X1 port map( G => n5110, D => n5005, Q => 
                           registers_9_26_port);
   registers_reg_9_25_inst : DLH_X1 port map( G => n5110, D => n5008, Q => 
                           registers_9_25_port);
   registers_reg_9_24_inst : DLH_X1 port map( G => n5110, D => n5011, Q => 
                           registers_9_24_port);
   registers_reg_9_23_inst : DLH_X1 port map( G => n5110, D => n5014, Q => 
                           registers_9_23_port);
   registers_reg_9_22_inst : DLH_X1 port map( G => n5110, D => n5017, Q => 
                           registers_9_22_port);
   registers_reg_9_21_inst : DLH_X1 port map( G => n5109, D => n5020, Q => 
                           registers_9_21_port);
   registers_reg_9_20_inst : DLH_X1 port map( G => n5109, D => n5023, Q => 
                           registers_9_20_port);
   registers_reg_9_19_inst : DLH_X1 port map( G => n5109, D => n5026, Q => 
                           registers_9_19_port);
   registers_reg_9_18_inst : DLH_X1 port map( G => n5109, D => n5029, Q => 
                           registers_9_18_port);
   registers_reg_9_17_inst : DLH_X1 port map( G => n5109, D => n5032, Q => 
                           registers_9_17_port);
   registers_reg_9_16_inst : DLH_X1 port map( G => n5109, D => n5035, Q => 
                           registers_9_16_port);
   registers_reg_9_15_inst : DLH_X1 port map( G => n5109, D => n5038, Q => 
                           registers_9_15_port);
   registers_reg_9_14_inst : DLH_X1 port map( G => n5109, D => n5041, Q => 
                           registers_9_14_port);
   registers_reg_9_13_inst : DLH_X1 port map( G => n5109, D => n5044, Q => 
                           registers_9_13_port);
   registers_reg_9_12_inst : DLH_X1 port map( G => n5109, D => n5047, Q => 
                           registers_9_12_port);
   registers_reg_9_11_inst : DLH_X1 port map( G => n5109, D => n5050, Q => 
                           registers_9_11_port);
   registers_reg_9_10_inst : DLH_X1 port map( G => n5108, D => n5053, Q => 
                           registers_9_10_port);
   registers_reg_9_9_inst : DLH_X1 port map( G => n5108, D => n5056, Q => 
                           registers_9_9_port);
   registers_reg_9_8_inst : DLH_X1 port map( G => n5108, D => n5059, Q => 
                           registers_9_8_port);
   registers_reg_9_7_inst : DLH_X1 port map( G => n5108, D => n5062, Q => 
                           registers_9_7_port);
   registers_reg_9_6_inst : DLH_X1 port map( G => n5108, D => n5065, Q => 
                           registers_9_6_port);
   registers_reg_9_5_inst : DLH_X1 port map( G => n5108, D => n5068, Q => 
                           registers_9_5_port);
   registers_reg_9_4_inst : DLH_X1 port map( G => n5108, D => n5071, Q => 
                           registers_9_4_port);
   registers_reg_9_3_inst : DLH_X1 port map( G => n5108, D => n5074, Q => 
                           registers_9_3_port);
   registers_reg_9_2_inst : DLH_X1 port map( G => n5108, D => n5077, Q => 
                           registers_9_2_port);
   registers_reg_9_1_inst : DLH_X1 port map( G => n5108, D => n5080, Q => 
                           registers_9_1_port);
   registers_reg_9_0_inst : DLH_X1 port map( G => n5108, D => n5083, Q => 
                           registers_9_0_port);
   registers_reg_10_31_inst : DLH_X1 port map( G => n5113, D => n4990, Q => 
                           registers_10_31_port);
   registers_reg_10_30_inst : DLH_X1 port map( G => n5113, D => n4993, Q => 
                           registers_10_30_port);
   registers_reg_10_29_inst : DLH_X1 port map( G => n5113, D => n4996, Q => 
                           registers_10_29_port);
   registers_reg_10_28_inst : DLH_X1 port map( G => n5113, D => n4999, Q => 
                           registers_10_28_port);
   registers_reg_10_27_inst : DLH_X1 port map( G => n5113, D => n5002, Q => 
                           registers_10_27_port);
   registers_reg_10_26_inst : DLH_X1 port map( G => n5113, D => n5005, Q => 
                           registers_10_26_port);
   registers_reg_10_25_inst : DLH_X1 port map( G => n5113, D => n5008, Q => 
                           registers_10_25_port);
   registers_reg_10_24_inst : DLH_X1 port map( G => n5113, D => n5011, Q => 
                           registers_10_24_port);
   registers_reg_10_23_inst : DLH_X1 port map( G => n5113, D => n5014, Q => 
                           registers_10_23_port);
   registers_reg_10_22_inst : DLH_X1 port map( G => n5113, D => n5017, Q => 
                           registers_10_22_port);
   registers_reg_10_21_inst : DLH_X1 port map( G => n5112, D => n5020, Q => 
                           registers_10_21_port);
   registers_reg_10_20_inst : DLH_X1 port map( G => n5112, D => n5023, Q => 
                           registers_10_20_port);
   registers_reg_10_19_inst : DLH_X1 port map( G => n5112, D => n5026, Q => 
                           registers_10_19_port);
   registers_reg_10_18_inst : DLH_X1 port map( G => n5112, D => n5029, Q => 
                           registers_10_18_port);
   registers_reg_10_17_inst : DLH_X1 port map( G => n5112, D => n5032, Q => 
                           registers_10_17_port);
   registers_reg_10_16_inst : DLH_X1 port map( G => n5112, D => n5035, Q => 
                           registers_10_16_port);
   registers_reg_10_15_inst : DLH_X1 port map( G => n5112, D => n5038, Q => 
                           registers_10_15_port);
   registers_reg_10_14_inst : DLH_X1 port map( G => n5112, D => n5041, Q => 
                           registers_10_14_port);
   registers_reg_10_13_inst : DLH_X1 port map( G => n5112, D => n5044, Q => 
                           registers_10_13_port);
   registers_reg_10_12_inst : DLH_X1 port map( G => n5112, D => n5047, Q => 
                           registers_10_12_port);
   registers_reg_10_11_inst : DLH_X1 port map( G => n5112, D => n5050, Q => 
                           registers_10_11_port);
   registers_reg_10_10_inst : DLH_X1 port map( G => n5111, D => n5053, Q => 
                           registers_10_10_port);
   registers_reg_10_9_inst : DLH_X1 port map( G => n5111, D => n5056, Q => 
                           registers_10_9_port);
   registers_reg_10_8_inst : DLH_X1 port map( G => n5111, D => n5059, Q => 
                           registers_10_8_port);
   registers_reg_10_7_inst : DLH_X1 port map( G => n5111, D => n5062, Q => 
                           registers_10_7_port);
   registers_reg_10_6_inst : DLH_X1 port map( G => n5111, D => n5065, Q => 
                           registers_10_6_port);
   registers_reg_10_5_inst : DLH_X1 port map( G => n5111, D => n5068, Q => 
                           registers_10_5_port);
   registers_reg_10_4_inst : DLH_X1 port map( G => n5111, D => n5071, Q => 
                           registers_10_4_port);
   registers_reg_10_3_inst : DLH_X1 port map( G => n5111, D => n5074, Q => 
                           registers_10_3_port);
   registers_reg_10_2_inst : DLH_X1 port map( G => n5111, D => n5077, Q => 
                           registers_10_2_port);
   registers_reg_10_1_inst : DLH_X1 port map( G => n5111, D => n5080, Q => 
                           registers_10_1_port);
   registers_reg_10_0_inst : DLH_X1 port map( G => n5111, D => n5083, Q => 
                           registers_10_0_port);
   registers_reg_11_31_inst : DLH_X1 port map( G => n5116, D => n4990, Q => 
                           registers_11_31_port);
   registers_reg_11_30_inst : DLH_X1 port map( G => n5116, D => n4993, Q => 
                           registers_11_30_port);
   registers_reg_11_29_inst : DLH_X1 port map( G => n5116, D => n4996, Q => 
                           registers_11_29_port);
   registers_reg_11_28_inst : DLH_X1 port map( G => n5116, D => n4999, Q => 
                           registers_11_28_port);
   registers_reg_11_27_inst : DLH_X1 port map( G => n5116, D => n5002, Q => 
                           registers_11_27_port);
   registers_reg_11_26_inst : DLH_X1 port map( G => n5116, D => n5005, Q => 
                           registers_11_26_port);
   registers_reg_11_25_inst : DLH_X1 port map( G => n5116, D => n5008, Q => 
                           registers_11_25_port);
   registers_reg_11_24_inst : DLH_X1 port map( G => n5116, D => n5011, Q => 
                           registers_11_24_port);
   registers_reg_11_23_inst : DLH_X1 port map( G => n5116, D => n5014, Q => 
                           registers_11_23_port);
   registers_reg_11_22_inst : DLH_X1 port map( G => n5116, D => n5017, Q => 
                           registers_11_22_port);
   registers_reg_11_21_inst : DLH_X1 port map( G => n5115, D => n5020, Q => 
                           registers_11_21_port);
   registers_reg_11_20_inst : DLH_X1 port map( G => n5115, D => n5023, Q => 
                           registers_11_20_port);
   registers_reg_11_19_inst : DLH_X1 port map( G => n5115, D => n5026, Q => 
                           registers_11_19_port);
   registers_reg_11_18_inst : DLH_X1 port map( G => n5115, D => n5029, Q => 
                           registers_11_18_port);
   registers_reg_11_17_inst : DLH_X1 port map( G => n5115, D => n5032, Q => 
                           registers_11_17_port);
   registers_reg_11_16_inst : DLH_X1 port map( G => n5115, D => n5035, Q => 
                           registers_11_16_port);
   registers_reg_11_15_inst : DLH_X1 port map( G => n5115, D => n5038, Q => 
                           registers_11_15_port);
   registers_reg_11_14_inst : DLH_X1 port map( G => n5115, D => n5041, Q => 
                           registers_11_14_port);
   registers_reg_11_13_inst : DLH_X1 port map( G => n5115, D => n5044, Q => 
                           registers_11_13_port);
   registers_reg_11_12_inst : DLH_X1 port map( G => n5115, D => n5047, Q => 
                           registers_11_12_port);
   registers_reg_11_11_inst : DLH_X1 port map( G => n5115, D => n5050, Q => 
                           registers_11_11_port);
   registers_reg_11_10_inst : DLH_X1 port map( G => n5114, D => n5053, Q => 
                           registers_11_10_port);
   registers_reg_11_9_inst : DLH_X1 port map( G => n5114, D => n5056, Q => 
                           registers_11_9_port);
   registers_reg_11_8_inst : DLH_X1 port map( G => n5114, D => n5059, Q => 
                           registers_11_8_port);
   registers_reg_11_7_inst : DLH_X1 port map( G => n5114, D => n5062, Q => 
                           registers_11_7_port);
   registers_reg_11_6_inst : DLH_X1 port map( G => n5114, D => n5065, Q => 
                           registers_11_6_port);
   registers_reg_11_5_inst : DLH_X1 port map( G => n5114, D => n5068, Q => 
                           registers_11_5_port);
   registers_reg_11_4_inst : DLH_X1 port map( G => n5114, D => n5071, Q => 
                           registers_11_4_port);
   registers_reg_11_3_inst : DLH_X1 port map( G => n5114, D => n5074, Q => 
                           registers_11_3_port);
   registers_reg_11_2_inst : DLH_X1 port map( G => n5114, D => n5077, Q => 
                           registers_11_2_port);
   registers_reg_11_1_inst : DLH_X1 port map( G => n5114, D => n5080, Q => 
                           registers_11_1_port);
   registers_reg_11_0_inst : DLH_X1 port map( G => n5114, D => n5083, Q => 
                           registers_11_0_port);
   registers_reg_12_31_inst : DLH_X1 port map( G => n5119, D => n4988, Q => 
                           registers_12_31_port);
   registers_reg_12_30_inst : DLH_X1 port map( G => n5119, D => n4991, Q => 
                           registers_12_30_port);
   registers_reg_12_29_inst : DLH_X1 port map( G => n5119, D => n4994, Q => 
                           registers_12_29_port);
   registers_reg_12_28_inst : DLH_X1 port map( G => n5119, D => n4997, Q => 
                           registers_12_28_port);
   registers_reg_12_27_inst : DLH_X1 port map( G => n5119, D => n5000, Q => 
                           registers_12_27_port);
   registers_reg_12_26_inst : DLH_X1 port map( G => n5119, D => n5003, Q => 
                           registers_12_26_port);
   registers_reg_12_25_inst : DLH_X1 port map( G => n5119, D => n5006, Q => 
                           registers_12_25_port);
   registers_reg_12_24_inst : DLH_X1 port map( G => n5119, D => n5009, Q => 
                           registers_12_24_port);
   registers_reg_12_23_inst : DLH_X1 port map( G => n5119, D => n5012, Q => 
                           registers_12_23_port);
   registers_reg_12_22_inst : DLH_X1 port map( G => n5119, D => n5015, Q => 
                           registers_12_22_port);
   registers_reg_12_21_inst : DLH_X1 port map( G => n5118, D => n5018, Q => 
                           registers_12_21_port);
   registers_reg_12_20_inst : DLH_X1 port map( G => n5118, D => n5021, Q => 
                           registers_12_20_port);
   registers_reg_12_19_inst : DLH_X1 port map( G => n5118, D => n5024, Q => 
                           registers_12_19_port);
   registers_reg_12_18_inst : DLH_X1 port map( G => n5118, D => n5027, Q => 
                           registers_12_18_port);
   registers_reg_12_17_inst : DLH_X1 port map( G => n5118, D => n5030, Q => 
                           registers_12_17_port);
   registers_reg_12_16_inst : DLH_X1 port map( G => n5118, D => n5033, Q => 
                           registers_12_16_port);
   registers_reg_12_15_inst : DLH_X1 port map( G => n5118, D => n5036, Q => 
                           registers_12_15_port);
   registers_reg_12_14_inst : DLH_X1 port map( G => n5118, D => n5039, Q => 
                           registers_12_14_port);
   registers_reg_12_13_inst : DLH_X1 port map( G => n5118, D => n5042, Q => 
                           registers_12_13_port);
   registers_reg_12_12_inst : DLH_X1 port map( G => n5118, D => n5045, Q => 
                           registers_12_12_port);
   registers_reg_12_11_inst : DLH_X1 port map( G => n5118, D => n5048, Q => 
                           registers_12_11_port);
   registers_reg_12_10_inst : DLH_X1 port map( G => n5117, D => n5051, Q => 
                           registers_12_10_port);
   registers_reg_12_9_inst : DLH_X1 port map( G => n5117, D => n5054, Q => 
                           registers_12_9_port);
   registers_reg_12_8_inst : DLH_X1 port map( G => n5117, D => n5057, Q => 
                           registers_12_8_port);
   registers_reg_12_7_inst : DLH_X1 port map( G => n5117, D => n5060, Q => 
                           registers_12_7_port);
   registers_reg_12_6_inst : DLH_X1 port map( G => n5117, D => n5063, Q => 
                           registers_12_6_port);
   registers_reg_12_5_inst : DLH_X1 port map( G => n5117, D => n5066, Q => 
                           registers_12_5_port);
   registers_reg_12_4_inst : DLH_X1 port map( G => n5117, D => n5069, Q => 
                           registers_12_4_port);
   registers_reg_12_3_inst : DLH_X1 port map( G => n5117, D => n5072, Q => 
                           registers_12_3_port);
   registers_reg_12_2_inst : DLH_X1 port map( G => n5117, D => n5075, Q => 
                           registers_12_2_port);
   registers_reg_12_1_inst : DLH_X1 port map( G => n5117, D => n5078, Q => 
                           registers_12_1_port);
   registers_reg_12_0_inst : DLH_X1 port map( G => n5117, D => n5081, Q => 
                           registers_12_0_port);
   registers_reg_13_31_inst : DLH_X1 port map( G => n5122, D => n4988, Q => 
                           registers_13_31_port);
   registers_reg_13_30_inst : DLH_X1 port map( G => n5122, D => n4991, Q => 
                           registers_13_30_port);
   registers_reg_13_29_inst : DLH_X1 port map( G => n5122, D => n4994, Q => 
                           registers_13_29_port);
   registers_reg_13_28_inst : DLH_X1 port map( G => n5122, D => n4997, Q => 
                           registers_13_28_port);
   registers_reg_13_27_inst : DLH_X1 port map( G => n5122, D => n5000, Q => 
                           registers_13_27_port);
   registers_reg_13_26_inst : DLH_X1 port map( G => n5122, D => n5003, Q => 
                           registers_13_26_port);
   registers_reg_13_25_inst : DLH_X1 port map( G => n5122, D => n5006, Q => 
                           registers_13_25_port);
   registers_reg_13_24_inst : DLH_X1 port map( G => n5122, D => n5009, Q => 
                           registers_13_24_port);
   registers_reg_13_23_inst : DLH_X1 port map( G => n5122, D => n5012, Q => 
                           registers_13_23_port);
   registers_reg_13_22_inst : DLH_X1 port map( G => n5122, D => n5015, Q => 
                           registers_13_22_port);
   registers_reg_13_21_inst : DLH_X1 port map( G => n5121, D => n5018, Q => 
                           registers_13_21_port);
   registers_reg_13_20_inst : DLH_X1 port map( G => n5121, D => n5021, Q => 
                           registers_13_20_port);
   registers_reg_13_19_inst : DLH_X1 port map( G => n5121, D => n5024, Q => 
                           registers_13_19_port);
   registers_reg_13_18_inst : DLH_X1 port map( G => n5121, D => n5027, Q => 
                           registers_13_18_port);
   registers_reg_13_17_inst : DLH_X1 port map( G => n5121, D => n5030, Q => 
                           registers_13_17_port);
   registers_reg_13_16_inst : DLH_X1 port map( G => n5121, D => n5033, Q => 
                           registers_13_16_port);
   registers_reg_13_15_inst : DLH_X1 port map( G => n5121, D => n5036, Q => 
                           registers_13_15_port);
   registers_reg_13_14_inst : DLH_X1 port map( G => n5121, D => n5039, Q => 
                           registers_13_14_port);
   registers_reg_13_13_inst : DLH_X1 port map( G => n5121, D => n5042, Q => 
                           registers_13_13_port);
   registers_reg_13_12_inst : DLH_X1 port map( G => n5121, D => n5045, Q => 
                           registers_13_12_port);
   registers_reg_13_11_inst : DLH_X1 port map( G => n5121, D => n5048, Q => 
                           registers_13_11_port);
   registers_reg_13_10_inst : DLH_X1 port map( G => n5120, D => n5051, Q => 
                           registers_13_10_port);
   registers_reg_13_9_inst : DLH_X1 port map( G => n5120, D => n5054, Q => 
                           registers_13_9_port);
   registers_reg_13_8_inst : DLH_X1 port map( G => n5120, D => n5057, Q => 
                           registers_13_8_port);
   registers_reg_13_7_inst : DLH_X1 port map( G => n5120, D => n5060, Q => 
                           registers_13_7_port);
   registers_reg_13_6_inst : DLH_X1 port map( G => n5120, D => n5063, Q => 
                           registers_13_6_port);
   registers_reg_13_5_inst : DLH_X1 port map( G => n5120, D => n5066, Q => 
                           registers_13_5_port);
   registers_reg_13_4_inst : DLH_X1 port map( G => n5120, D => n5069, Q => 
                           registers_13_4_port);
   registers_reg_13_3_inst : DLH_X1 port map( G => n5120, D => n5072, Q => 
                           registers_13_3_port);
   registers_reg_13_2_inst : DLH_X1 port map( G => n5120, D => n5075, Q => 
                           registers_13_2_port);
   registers_reg_13_1_inst : DLH_X1 port map( G => n5120, D => n5078, Q => 
                           registers_13_1_port);
   registers_reg_13_0_inst : DLH_X1 port map( G => n5120, D => n5081, Q => 
                           registers_13_0_port);
   registers_reg_14_31_inst : DLH_X1 port map( G => n5125, D => n4988, Q => 
                           registers_14_31_port);
   registers_reg_14_30_inst : DLH_X1 port map( G => n5125, D => n4991, Q => 
                           registers_14_30_port);
   registers_reg_14_29_inst : DLH_X1 port map( G => n5125, D => n4994, Q => 
                           registers_14_29_port);
   registers_reg_14_28_inst : DLH_X1 port map( G => n5125, D => n4997, Q => 
                           registers_14_28_port);
   registers_reg_14_27_inst : DLH_X1 port map( G => n5125, D => n5000, Q => 
                           registers_14_27_port);
   registers_reg_14_26_inst : DLH_X1 port map( G => n5125, D => n5003, Q => 
                           registers_14_26_port);
   registers_reg_14_25_inst : DLH_X1 port map( G => n5125, D => n5006, Q => 
                           registers_14_25_port);
   registers_reg_14_24_inst : DLH_X1 port map( G => n5125, D => n5009, Q => 
                           registers_14_24_port);
   registers_reg_14_23_inst : DLH_X1 port map( G => n5125, D => n5012, Q => 
                           registers_14_23_port);
   registers_reg_14_22_inst : DLH_X1 port map( G => n5125, D => n5015, Q => 
                           registers_14_22_port);
   registers_reg_14_21_inst : DLH_X1 port map( G => n5124, D => n5018, Q => 
                           registers_14_21_port);
   registers_reg_14_20_inst : DLH_X1 port map( G => n5124, D => n5021, Q => 
                           registers_14_20_port);
   registers_reg_14_19_inst : DLH_X1 port map( G => n5124, D => n5024, Q => 
                           registers_14_19_port);
   registers_reg_14_18_inst : DLH_X1 port map( G => n5124, D => n5027, Q => 
                           registers_14_18_port);
   registers_reg_14_17_inst : DLH_X1 port map( G => n5124, D => n5030, Q => 
                           registers_14_17_port);
   registers_reg_14_16_inst : DLH_X1 port map( G => n5124, D => n5033, Q => 
                           registers_14_16_port);
   registers_reg_14_15_inst : DLH_X1 port map( G => n5124, D => n5036, Q => 
                           registers_14_15_port);
   registers_reg_14_14_inst : DLH_X1 port map( G => n5124, D => n5039, Q => 
                           registers_14_14_port);
   registers_reg_14_13_inst : DLH_X1 port map( G => n5124, D => n5042, Q => 
                           registers_14_13_port);
   registers_reg_14_12_inst : DLH_X1 port map( G => n5124, D => n5045, Q => 
                           registers_14_12_port);
   registers_reg_14_11_inst : DLH_X1 port map( G => n5124, D => n5048, Q => 
                           registers_14_11_port);
   registers_reg_14_10_inst : DLH_X1 port map( G => n5123, D => n5051, Q => 
                           registers_14_10_port);
   registers_reg_14_9_inst : DLH_X1 port map( G => n5123, D => n5054, Q => 
                           registers_14_9_port);
   registers_reg_14_8_inst : DLH_X1 port map( G => n5123, D => n5057, Q => 
                           registers_14_8_port);
   registers_reg_14_7_inst : DLH_X1 port map( G => n5123, D => n5060, Q => 
                           registers_14_7_port);
   registers_reg_14_6_inst : DLH_X1 port map( G => n5123, D => n5063, Q => 
                           registers_14_6_port);
   registers_reg_14_5_inst : DLH_X1 port map( G => n5123, D => n5066, Q => 
                           registers_14_5_port);
   registers_reg_14_4_inst : DLH_X1 port map( G => n5123, D => n5069, Q => 
                           registers_14_4_port);
   registers_reg_14_3_inst : DLH_X1 port map( G => n5123, D => n5072, Q => 
                           registers_14_3_port);
   registers_reg_14_2_inst : DLH_X1 port map( G => n5123, D => n5075, Q => 
                           registers_14_2_port);
   registers_reg_14_1_inst : DLH_X1 port map( G => n5123, D => n5078, Q => 
                           registers_14_1_port);
   registers_reg_14_0_inst : DLH_X1 port map( G => n5123, D => n5081, Q => 
                           registers_14_0_port);
   registers_reg_15_31_inst : DLH_X1 port map( G => n5128, D => n4988, Q => 
                           registers_15_31_port);
   registers_reg_15_30_inst : DLH_X1 port map( G => n5128, D => n4991, Q => 
                           registers_15_30_port);
   registers_reg_15_29_inst : DLH_X1 port map( G => n5128, D => n4994, Q => 
                           registers_15_29_port);
   registers_reg_15_28_inst : DLH_X1 port map( G => n5128, D => n4997, Q => 
                           registers_15_28_port);
   registers_reg_15_27_inst : DLH_X1 port map( G => n5128, D => n5000, Q => 
                           registers_15_27_port);
   registers_reg_15_26_inst : DLH_X1 port map( G => n5128, D => n5003, Q => 
                           registers_15_26_port);
   registers_reg_15_25_inst : DLH_X1 port map( G => n5128, D => n5006, Q => 
                           registers_15_25_port);
   registers_reg_15_24_inst : DLH_X1 port map( G => n5128, D => n5009, Q => 
                           registers_15_24_port);
   registers_reg_15_23_inst : DLH_X1 port map( G => n5128, D => n5012, Q => 
                           registers_15_23_port);
   registers_reg_15_22_inst : DLH_X1 port map( G => n5128, D => n5015, Q => 
                           registers_15_22_port);
   registers_reg_15_21_inst : DLH_X1 port map( G => n5127, D => n5018, Q => 
                           registers_15_21_port);
   registers_reg_15_20_inst : DLH_X1 port map( G => n5127, D => n5021, Q => 
                           registers_15_20_port);
   registers_reg_15_19_inst : DLH_X1 port map( G => n5127, D => n5024, Q => 
                           registers_15_19_port);
   registers_reg_15_18_inst : DLH_X1 port map( G => n5127, D => n5027, Q => 
                           registers_15_18_port);
   registers_reg_15_17_inst : DLH_X1 port map( G => n5127, D => n5030, Q => 
                           registers_15_17_port);
   registers_reg_15_16_inst : DLH_X1 port map( G => n5127, D => n5033, Q => 
                           registers_15_16_port);
   registers_reg_15_15_inst : DLH_X1 port map( G => n5127, D => n5036, Q => 
                           registers_15_15_port);
   registers_reg_15_14_inst : DLH_X1 port map( G => n5127, D => n5039, Q => 
                           registers_15_14_port);
   registers_reg_15_13_inst : DLH_X1 port map( G => n5127, D => n5042, Q => 
                           registers_15_13_port);
   registers_reg_15_12_inst : DLH_X1 port map( G => n5127, D => n5045, Q => 
                           registers_15_12_port);
   registers_reg_15_11_inst : DLH_X1 port map( G => n5127, D => n5048, Q => 
                           registers_15_11_port);
   registers_reg_15_10_inst : DLH_X1 port map( G => n5126, D => n5051, Q => 
                           registers_15_10_port);
   registers_reg_15_9_inst : DLH_X1 port map( G => n5126, D => n5054, Q => 
                           registers_15_9_port);
   registers_reg_15_8_inst : DLH_X1 port map( G => n5126, D => n5057, Q => 
                           registers_15_8_port);
   registers_reg_15_7_inst : DLH_X1 port map( G => n5126, D => n5060, Q => 
                           registers_15_7_port);
   registers_reg_15_6_inst : DLH_X1 port map( G => n5126, D => n5063, Q => 
                           registers_15_6_port);
   registers_reg_15_5_inst : DLH_X1 port map( G => n5126, D => n5066, Q => 
                           registers_15_5_port);
   registers_reg_15_4_inst : DLH_X1 port map( G => n5126, D => n5069, Q => 
                           registers_15_4_port);
   registers_reg_15_3_inst : DLH_X1 port map( G => n5126, D => n5072, Q => 
                           registers_15_3_port);
   registers_reg_15_2_inst : DLH_X1 port map( G => n5126, D => n5075, Q => 
                           registers_15_2_port);
   registers_reg_15_1_inst : DLH_X1 port map( G => n5126, D => n5078, Q => 
                           registers_15_1_port);
   registers_reg_15_0_inst : DLH_X1 port map( G => n5126, D => n5081, Q => 
                           registers_15_0_port);
   registers_reg_16_31_inst : DLH_X1 port map( G => n5131, D => n4988, Q => 
                           registers_16_31_port);
   registers_reg_16_30_inst : DLH_X1 port map( G => n5131, D => n4991, Q => 
                           registers_16_30_port);
   registers_reg_16_29_inst : DLH_X1 port map( G => n5131, D => n4994, Q => 
                           registers_16_29_port);
   registers_reg_16_28_inst : DLH_X1 port map( G => n5131, D => n4997, Q => 
                           registers_16_28_port);
   registers_reg_16_27_inst : DLH_X1 port map( G => n5131, D => n5000, Q => 
                           registers_16_27_port);
   registers_reg_16_26_inst : DLH_X1 port map( G => n5131, D => n5003, Q => 
                           registers_16_26_port);
   registers_reg_16_25_inst : DLH_X1 port map( G => n5131, D => n5006, Q => 
                           registers_16_25_port);
   registers_reg_16_24_inst : DLH_X1 port map( G => n5131, D => n5009, Q => 
                           registers_16_24_port);
   registers_reg_16_23_inst : DLH_X1 port map( G => n5131, D => n5012, Q => 
                           registers_16_23_port);
   registers_reg_16_22_inst : DLH_X1 port map( G => n5131, D => n5015, Q => 
                           registers_16_22_port);
   registers_reg_16_21_inst : DLH_X1 port map( G => n5130, D => n5018, Q => 
                           registers_16_21_port);
   registers_reg_16_20_inst : DLH_X1 port map( G => n5130, D => n5021, Q => 
                           registers_16_20_port);
   registers_reg_16_19_inst : DLH_X1 port map( G => n5130, D => n5024, Q => 
                           registers_16_19_port);
   registers_reg_16_18_inst : DLH_X1 port map( G => n5130, D => n5027, Q => 
                           registers_16_18_port);
   registers_reg_16_17_inst : DLH_X1 port map( G => n5130, D => n5030, Q => 
                           registers_16_17_port);
   registers_reg_16_16_inst : DLH_X1 port map( G => n5130, D => n5033, Q => 
                           registers_16_16_port);
   registers_reg_16_15_inst : DLH_X1 port map( G => n5130, D => n5036, Q => 
                           registers_16_15_port);
   registers_reg_16_14_inst : DLH_X1 port map( G => n5130, D => n5039, Q => 
                           registers_16_14_port);
   registers_reg_16_13_inst : DLH_X1 port map( G => n5130, D => n5042, Q => 
                           registers_16_13_port);
   registers_reg_16_12_inst : DLH_X1 port map( G => n5130, D => n5045, Q => 
                           registers_16_12_port);
   registers_reg_16_11_inst : DLH_X1 port map( G => n5130, D => n5048, Q => 
                           registers_16_11_port);
   registers_reg_16_10_inst : DLH_X1 port map( G => n5129, D => n5051, Q => 
                           registers_16_10_port);
   registers_reg_16_9_inst : DLH_X1 port map( G => n5129, D => n5054, Q => 
                           registers_16_9_port);
   registers_reg_16_8_inst : DLH_X1 port map( G => n5129, D => n5057, Q => 
                           registers_16_8_port);
   registers_reg_16_7_inst : DLH_X1 port map( G => n5129, D => n5060, Q => 
                           registers_16_7_port);
   registers_reg_16_6_inst : DLH_X1 port map( G => n5129, D => n5063, Q => 
                           registers_16_6_port);
   registers_reg_16_5_inst : DLH_X1 port map( G => n5129, D => n5066, Q => 
                           registers_16_5_port);
   registers_reg_16_4_inst : DLH_X1 port map( G => n5129, D => n5069, Q => 
                           registers_16_4_port);
   registers_reg_16_3_inst : DLH_X1 port map( G => n5129, D => n5072, Q => 
                           registers_16_3_port);
   registers_reg_16_2_inst : DLH_X1 port map( G => n5129, D => n5075, Q => 
                           registers_16_2_port);
   registers_reg_16_1_inst : DLH_X1 port map( G => n5129, D => n5078, Q => 
                           registers_16_1_port);
   registers_reg_16_0_inst : DLH_X1 port map( G => n5129, D => n5081, Q => 
                           registers_16_0_port);
   registers_reg_17_31_inst : DLH_X1 port map( G => n5134, D => n4988, Q => 
                           registers_17_31_port);
   registers_reg_17_30_inst : DLH_X1 port map( G => n5134, D => n4991, Q => 
                           registers_17_30_port);
   registers_reg_17_29_inst : DLH_X1 port map( G => n5134, D => n4994, Q => 
                           registers_17_29_port);
   registers_reg_17_28_inst : DLH_X1 port map( G => n5134, D => n4997, Q => 
                           registers_17_28_port);
   registers_reg_17_27_inst : DLH_X1 port map( G => n5134, D => n5000, Q => 
                           registers_17_27_port);
   registers_reg_17_26_inst : DLH_X1 port map( G => n5134, D => n5003, Q => 
                           registers_17_26_port);
   registers_reg_17_25_inst : DLH_X1 port map( G => n5134, D => n5006, Q => 
                           registers_17_25_port);
   registers_reg_17_24_inst : DLH_X1 port map( G => n5134, D => n5009, Q => 
                           registers_17_24_port);
   registers_reg_17_23_inst : DLH_X1 port map( G => n5134, D => n5012, Q => 
                           registers_17_23_port);
   registers_reg_17_22_inst : DLH_X1 port map( G => n5134, D => n5015, Q => 
                           registers_17_22_port);
   registers_reg_17_21_inst : DLH_X1 port map( G => n5133, D => n5018, Q => 
                           registers_17_21_port);
   registers_reg_17_20_inst : DLH_X1 port map( G => n5133, D => n5021, Q => 
                           registers_17_20_port);
   registers_reg_17_19_inst : DLH_X1 port map( G => n5133, D => n5024, Q => 
                           registers_17_19_port);
   registers_reg_17_18_inst : DLH_X1 port map( G => n5133, D => n5027, Q => 
                           registers_17_18_port);
   registers_reg_17_17_inst : DLH_X1 port map( G => n5133, D => n5030, Q => 
                           registers_17_17_port);
   registers_reg_17_16_inst : DLH_X1 port map( G => n5133, D => n5033, Q => 
                           registers_17_16_port);
   registers_reg_17_15_inst : DLH_X1 port map( G => n5133, D => n5036, Q => 
                           registers_17_15_port);
   registers_reg_17_14_inst : DLH_X1 port map( G => n5133, D => n5039, Q => 
                           registers_17_14_port);
   registers_reg_17_13_inst : DLH_X1 port map( G => n5133, D => n5042, Q => 
                           registers_17_13_port);
   registers_reg_17_12_inst : DLH_X1 port map( G => n5133, D => n5045, Q => 
                           registers_17_12_port);
   registers_reg_17_11_inst : DLH_X1 port map( G => n5133, D => n5048, Q => 
                           registers_17_11_port);
   registers_reg_17_10_inst : DLH_X1 port map( G => n5132, D => n5051, Q => 
                           registers_17_10_port);
   registers_reg_17_9_inst : DLH_X1 port map( G => n5132, D => n5054, Q => 
                           registers_17_9_port);
   registers_reg_17_8_inst : DLH_X1 port map( G => n5132, D => n5057, Q => 
                           registers_17_8_port);
   registers_reg_17_7_inst : DLH_X1 port map( G => n5132, D => n5060, Q => 
                           registers_17_7_port);
   registers_reg_17_6_inst : DLH_X1 port map( G => n5132, D => n5063, Q => 
                           registers_17_6_port);
   registers_reg_17_5_inst : DLH_X1 port map( G => n5132, D => n5066, Q => 
                           registers_17_5_port);
   registers_reg_17_4_inst : DLH_X1 port map( G => n5132, D => n5069, Q => 
                           registers_17_4_port);
   registers_reg_17_3_inst : DLH_X1 port map( G => n5132, D => n5072, Q => 
                           registers_17_3_port);
   registers_reg_17_2_inst : DLH_X1 port map( G => n5132, D => n5075, Q => 
                           registers_17_2_port);
   registers_reg_17_1_inst : DLH_X1 port map( G => n5132, D => n5078, Q => 
                           registers_17_1_port);
   registers_reg_17_0_inst : DLH_X1 port map( G => n5132, D => n5081, Q => 
                           registers_17_0_port);
   registers_reg_18_31_inst : DLH_X1 port map( G => n5137, D => n4988, Q => 
                           registers_18_31_port);
   registers_reg_18_30_inst : DLH_X1 port map( G => n5137, D => n4991, Q => 
                           registers_18_30_port);
   registers_reg_18_29_inst : DLH_X1 port map( G => n5137, D => n4994, Q => 
                           registers_18_29_port);
   registers_reg_18_28_inst : DLH_X1 port map( G => n5137, D => n4997, Q => 
                           registers_18_28_port);
   registers_reg_18_27_inst : DLH_X1 port map( G => n5137, D => n5000, Q => 
                           registers_18_27_port);
   registers_reg_18_26_inst : DLH_X1 port map( G => n5137, D => n5003, Q => 
                           registers_18_26_port);
   registers_reg_18_25_inst : DLH_X1 port map( G => n5137, D => n5006, Q => 
                           registers_18_25_port);
   registers_reg_18_24_inst : DLH_X1 port map( G => n5137, D => n5009, Q => 
                           registers_18_24_port);
   registers_reg_18_23_inst : DLH_X1 port map( G => n5137, D => n5012, Q => 
                           registers_18_23_port);
   registers_reg_18_22_inst : DLH_X1 port map( G => n5137, D => n5015, Q => 
                           registers_18_22_port);
   registers_reg_18_21_inst : DLH_X1 port map( G => n5136, D => n5018, Q => 
                           registers_18_21_port);
   registers_reg_18_20_inst : DLH_X1 port map( G => n5136, D => n5021, Q => 
                           registers_18_20_port);
   registers_reg_18_19_inst : DLH_X1 port map( G => n5136, D => n5024, Q => 
                           registers_18_19_port);
   registers_reg_18_18_inst : DLH_X1 port map( G => n5136, D => n5027, Q => 
                           registers_18_18_port);
   registers_reg_18_17_inst : DLH_X1 port map( G => n5136, D => n5030, Q => 
                           registers_18_17_port);
   registers_reg_18_16_inst : DLH_X1 port map( G => n5136, D => n5033, Q => 
                           registers_18_16_port);
   registers_reg_18_15_inst : DLH_X1 port map( G => n5136, D => n5036, Q => 
                           registers_18_15_port);
   registers_reg_18_14_inst : DLH_X1 port map( G => n5136, D => n5039, Q => 
                           registers_18_14_port);
   registers_reg_18_13_inst : DLH_X1 port map( G => n5136, D => n5042, Q => 
                           registers_18_13_port);
   registers_reg_18_12_inst : DLH_X1 port map( G => n5136, D => n5045, Q => 
                           registers_18_12_port);
   registers_reg_18_11_inst : DLH_X1 port map( G => n5136, D => n5048, Q => 
                           registers_18_11_port);
   registers_reg_18_10_inst : DLH_X1 port map( G => n5135, D => n5051, Q => 
                           registers_18_10_port);
   registers_reg_18_9_inst : DLH_X1 port map( G => n5135, D => n5054, Q => 
                           registers_18_9_port);
   registers_reg_18_8_inst : DLH_X1 port map( G => n5135, D => n5057, Q => 
                           registers_18_8_port);
   registers_reg_18_7_inst : DLH_X1 port map( G => n5135, D => n5060, Q => 
                           registers_18_7_port);
   registers_reg_18_6_inst : DLH_X1 port map( G => n5135, D => n5063, Q => 
                           registers_18_6_port);
   registers_reg_18_5_inst : DLH_X1 port map( G => n5135, D => n5066, Q => 
                           registers_18_5_port);
   registers_reg_18_4_inst : DLH_X1 port map( G => n5135, D => n5069, Q => 
                           registers_18_4_port);
   registers_reg_18_3_inst : DLH_X1 port map( G => n5135, D => n5072, Q => 
                           registers_18_3_port);
   registers_reg_18_2_inst : DLH_X1 port map( G => n5135, D => n5075, Q => 
                           registers_18_2_port);
   registers_reg_18_1_inst : DLH_X1 port map( G => n5135, D => n5078, Q => 
                           registers_18_1_port);
   registers_reg_18_0_inst : DLH_X1 port map( G => n5135, D => n5081, Q => 
                           registers_18_0_port);
   registers_reg_19_31_inst : DLH_X1 port map( G => n5140, D => n4988, Q => 
                           registers_19_31_port);
   registers_reg_19_30_inst : DLH_X1 port map( G => n5140, D => n4991, Q => 
                           registers_19_30_port);
   registers_reg_19_29_inst : DLH_X1 port map( G => n5140, D => n4994, Q => 
                           registers_19_29_port);
   registers_reg_19_28_inst : DLH_X1 port map( G => n5140, D => n4997, Q => 
                           registers_19_28_port);
   registers_reg_19_27_inst : DLH_X1 port map( G => n5140, D => n5000, Q => 
                           registers_19_27_port);
   registers_reg_19_26_inst : DLH_X1 port map( G => n5140, D => n5003, Q => 
                           registers_19_26_port);
   registers_reg_19_25_inst : DLH_X1 port map( G => n5140, D => n5006, Q => 
                           registers_19_25_port);
   registers_reg_19_24_inst : DLH_X1 port map( G => n5140, D => n5009, Q => 
                           registers_19_24_port);
   registers_reg_19_23_inst : DLH_X1 port map( G => n5140, D => n5012, Q => 
                           registers_19_23_port);
   registers_reg_19_22_inst : DLH_X1 port map( G => n5140, D => n5015, Q => 
                           registers_19_22_port);
   registers_reg_19_21_inst : DLH_X1 port map( G => n5139, D => n5018, Q => 
                           registers_19_21_port);
   registers_reg_19_20_inst : DLH_X1 port map( G => n5139, D => n5021, Q => 
                           registers_19_20_port);
   registers_reg_19_19_inst : DLH_X1 port map( G => n5139, D => n5024, Q => 
                           registers_19_19_port);
   registers_reg_19_18_inst : DLH_X1 port map( G => n5139, D => n5027, Q => 
                           registers_19_18_port);
   registers_reg_19_17_inst : DLH_X1 port map( G => n5139, D => n5030, Q => 
                           registers_19_17_port);
   registers_reg_19_16_inst : DLH_X1 port map( G => n5139, D => n5033, Q => 
                           registers_19_16_port);
   registers_reg_19_15_inst : DLH_X1 port map( G => n5139, D => n5036, Q => 
                           registers_19_15_port);
   registers_reg_19_14_inst : DLH_X1 port map( G => n5139, D => n5039, Q => 
                           registers_19_14_port);
   registers_reg_19_13_inst : DLH_X1 port map( G => n5139, D => n5042, Q => 
                           registers_19_13_port);
   registers_reg_19_12_inst : DLH_X1 port map( G => n5139, D => n5045, Q => 
                           registers_19_12_port);
   registers_reg_19_11_inst : DLH_X1 port map( G => n5139, D => n5048, Q => 
                           registers_19_11_port);
   registers_reg_19_10_inst : DLH_X1 port map( G => n5138, D => n5051, Q => 
                           registers_19_10_port);
   registers_reg_19_9_inst : DLH_X1 port map( G => n5138, D => n5054, Q => 
                           registers_19_9_port);
   registers_reg_19_8_inst : DLH_X1 port map( G => n5138, D => n5057, Q => 
                           registers_19_8_port);
   registers_reg_19_7_inst : DLH_X1 port map( G => n5138, D => n5060, Q => 
                           registers_19_7_port);
   registers_reg_19_6_inst : DLH_X1 port map( G => n5138, D => n5063, Q => 
                           registers_19_6_port);
   registers_reg_19_5_inst : DLH_X1 port map( G => n5138, D => n5066, Q => 
                           registers_19_5_port);
   registers_reg_19_4_inst : DLH_X1 port map( G => n5138, D => n5069, Q => 
                           registers_19_4_port);
   registers_reg_19_3_inst : DLH_X1 port map( G => n5138, D => n5072, Q => 
                           registers_19_3_port);
   registers_reg_19_2_inst : DLH_X1 port map( G => n5138, D => n5075, Q => 
                           registers_19_2_port);
   registers_reg_19_1_inst : DLH_X1 port map( G => n5138, D => n5078, Q => 
                           registers_19_1_port);
   registers_reg_19_0_inst : DLH_X1 port map( G => n5138, D => n5081, Q => 
                           registers_19_0_port);
   registers_reg_20_31_inst : DLH_X1 port map( G => n5143, D => n4988, Q => 
                           registers_20_31_port);
   registers_reg_20_30_inst : DLH_X1 port map( G => n5143, D => n4991, Q => 
                           registers_20_30_port);
   registers_reg_20_29_inst : DLH_X1 port map( G => n5143, D => n4994, Q => 
                           registers_20_29_port);
   registers_reg_20_28_inst : DLH_X1 port map( G => n5143, D => n4997, Q => 
                           registers_20_28_port);
   registers_reg_20_27_inst : DLH_X1 port map( G => n5143, D => n5000, Q => 
                           registers_20_27_port);
   registers_reg_20_26_inst : DLH_X1 port map( G => n5143, D => n5003, Q => 
                           registers_20_26_port);
   registers_reg_20_25_inst : DLH_X1 port map( G => n5143, D => n5006, Q => 
                           registers_20_25_port);
   registers_reg_20_24_inst : DLH_X1 port map( G => n5143, D => n5009, Q => 
                           registers_20_24_port);
   registers_reg_20_23_inst : DLH_X1 port map( G => n5143, D => n5012, Q => 
                           registers_20_23_port);
   registers_reg_20_22_inst : DLH_X1 port map( G => n5143, D => n5015, Q => 
                           registers_20_22_port);
   registers_reg_20_21_inst : DLH_X1 port map( G => n5142, D => n5018, Q => 
                           registers_20_21_port);
   registers_reg_20_20_inst : DLH_X1 port map( G => n5142, D => n5021, Q => 
                           registers_20_20_port);
   registers_reg_20_19_inst : DLH_X1 port map( G => n5142, D => n5024, Q => 
                           registers_20_19_port);
   registers_reg_20_18_inst : DLH_X1 port map( G => n5142, D => n5027, Q => 
                           registers_20_18_port);
   registers_reg_20_17_inst : DLH_X1 port map( G => n5142, D => n5030, Q => 
                           registers_20_17_port);
   registers_reg_20_16_inst : DLH_X1 port map( G => n5142, D => n5033, Q => 
                           registers_20_16_port);
   registers_reg_20_15_inst : DLH_X1 port map( G => n5142, D => n5036, Q => 
                           registers_20_15_port);
   registers_reg_20_14_inst : DLH_X1 port map( G => n5142, D => n5039, Q => 
                           registers_20_14_port);
   registers_reg_20_13_inst : DLH_X1 port map( G => n5142, D => n5042, Q => 
                           registers_20_13_port);
   registers_reg_20_12_inst : DLH_X1 port map( G => n5142, D => n5045, Q => 
                           registers_20_12_port);
   registers_reg_20_11_inst : DLH_X1 port map( G => n5142, D => n5048, Q => 
                           registers_20_11_port);
   registers_reg_20_10_inst : DLH_X1 port map( G => n5141, D => n5051, Q => 
                           registers_20_10_port);
   registers_reg_20_9_inst : DLH_X1 port map( G => n5141, D => n5054, Q => 
                           registers_20_9_port);
   registers_reg_20_8_inst : DLH_X1 port map( G => n5141, D => n5057, Q => 
                           registers_20_8_port);
   registers_reg_20_7_inst : DLH_X1 port map( G => n5141, D => n5060, Q => 
                           registers_20_7_port);
   registers_reg_20_6_inst : DLH_X1 port map( G => n5141, D => n5063, Q => 
                           registers_20_6_port);
   registers_reg_20_5_inst : DLH_X1 port map( G => n5141, D => n5066, Q => 
                           registers_20_5_port);
   registers_reg_20_4_inst : DLH_X1 port map( G => n5141, D => n5069, Q => 
                           registers_20_4_port);
   registers_reg_20_3_inst : DLH_X1 port map( G => n5141, D => n5072, Q => 
                           registers_20_3_port);
   registers_reg_20_2_inst : DLH_X1 port map( G => n5141, D => n5075, Q => 
                           registers_20_2_port);
   registers_reg_20_1_inst : DLH_X1 port map( G => n5141, D => n5078, Q => 
                           registers_20_1_port);
   registers_reg_20_0_inst : DLH_X1 port map( G => n5141, D => n5081, Q => 
                           registers_20_0_port);
   registers_reg_21_31_inst : DLH_X1 port map( G => n5146, D => n4989, Q => 
                           registers_21_31_port);
   registers_reg_21_30_inst : DLH_X1 port map( G => n5146, D => n4992, Q => 
                           registers_21_30_port);
   registers_reg_21_29_inst : DLH_X1 port map( G => n5146, D => n4995, Q => 
                           registers_21_29_port);
   registers_reg_21_28_inst : DLH_X1 port map( G => n5146, D => n4998, Q => 
                           registers_21_28_port);
   registers_reg_21_27_inst : DLH_X1 port map( G => n5146, D => n5001, Q => 
                           registers_21_27_port);
   registers_reg_21_26_inst : DLH_X1 port map( G => n5146, D => n5004, Q => 
                           registers_21_26_port);
   registers_reg_21_25_inst : DLH_X1 port map( G => n5146, D => n5007, Q => 
                           registers_21_25_port);
   registers_reg_21_24_inst : DLH_X1 port map( G => n5146, D => n5010, Q => 
                           registers_21_24_port);
   registers_reg_21_23_inst : DLH_X1 port map( G => n5146, D => n5013, Q => 
                           registers_21_23_port);
   registers_reg_21_22_inst : DLH_X1 port map( G => n5146, D => n5016, Q => 
                           registers_21_22_port);
   registers_reg_21_21_inst : DLH_X1 port map( G => n5145, D => n5019, Q => 
                           registers_21_21_port);
   registers_reg_21_20_inst : DLH_X1 port map( G => n5145, D => n5022, Q => 
                           registers_21_20_port);
   registers_reg_21_19_inst : DLH_X1 port map( G => n5145, D => n5025, Q => 
                           registers_21_19_port);
   registers_reg_21_18_inst : DLH_X1 port map( G => n5145, D => n5028, Q => 
                           registers_21_18_port);
   registers_reg_21_17_inst : DLH_X1 port map( G => n5145, D => n5031, Q => 
                           registers_21_17_port);
   registers_reg_21_16_inst : DLH_X1 port map( G => n5145, D => n5034, Q => 
                           registers_21_16_port);
   registers_reg_21_15_inst : DLH_X1 port map( G => n5145, D => n5037, Q => 
                           registers_21_15_port);
   registers_reg_21_14_inst : DLH_X1 port map( G => n5145, D => n5040, Q => 
                           registers_21_14_port);
   registers_reg_21_13_inst : DLH_X1 port map( G => n5145, D => n5043, Q => 
                           registers_21_13_port);
   registers_reg_21_12_inst : DLH_X1 port map( G => n5145, D => n5046, Q => 
                           registers_21_12_port);
   registers_reg_21_11_inst : DLH_X1 port map( G => n5145, D => n5049, Q => 
                           registers_21_11_port);
   registers_reg_21_10_inst : DLH_X1 port map( G => n5144, D => n5052, Q => 
                           registers_21_10_port);
   registers_reg_21_9_inst : DLH_X1 port map( G => n5144, D => n5055, Q => 
                           registers_21_9_port);
   registers_reg_21_8_inst : DLH_X1 port map( G => n5144, D => n5058, Q => 
                           registers_21_8_port);
   registers_reg_21_7_inst : DLH_X1 port map( G => n5144, D => n5061, Q => 
                           registers_21_7_port);
   registers_reg_21_6_inst : DLH_X1 port map( G => n5144, D => n5064, Q => 
                           registers_21_6_port);
   registers_reg_21_5_inst : DLH_X1 port map( G => n5144, D => n5067, Q => 
                           registers_21_5_port);
   registers_reg_21_4_inst : DLH_X1 port map( G => n5144, D => n5070, Q => 
                           registers_21_4_port);
   registers_reg_21_3_inst : DLH_X1 port map( G => n5144, D => n5073, Q => 
                           registers_21_3_port);
   registers_reg_21_2_inst : DLH_X1 port map( G => n5144, D => n5076, Q => 
                           registers_21_2_port);
   registers_reg_21_1_inst : DLH_X1 port map( G => n5144, D => n5079, Q => 
                           registers_21_1_port);
   registers_reg_21_0_inst : DLH_X1 port map( G => n5144, D => n5082, Q => 
                           registers_21_0_port);
   registers_reg_22_31_inst : DLH_X1 port map( G => n5149, D => n4989, Q => 
                           registers_22_31_port);
   registers_reg_22_30_inst : DLH_X1 port map( G => n5149, D => n4992, Q => 
                           registers_22_30_port);
   registers_reg_22_29_inst : DLH_X1 port map( G => n5149, D => n4995, Q => 
                           registers_22_29_port);
   registers_reg_22_28_inst : DLH_X1 port map( G => n5149, D => n4998, Q => 
                           registers_22_28_port);
   registers_reg_22_27_inst : DLH_X1 port map( G => n5149, D => n5001, Q => 
                           registers_22_27_port);
   registers_reg_22_26_inst : DLH_X1 port map( G => n5149, D => n5004, Q => 
                           registers_22_26_port);
   registers_reg_22_25_inst : DLH_X1 port map( G => n5149, D => n5007, Q => 
                           registers_22_25_port);
   registers_reg_22_24_inst : DLH_X1 port map( G => n5149, D => n5010, Q => 
                           registers_22_24_port);
   registers_reg_22_23_inst : DLH_X1 port map( G => n5149, D => n5013, Q => 
                           registers_22_23_port);
   registers_reg_22_22_inst : DLH_X1 port map( G => n5149, D => n5016, Q => 
                           registers_22_22_port);
   registers_reg_22_21_inst : DLH_X1 port map( G => n5148, D => n5019, Q => 
                           registers_22_21_port);
   registers_reg_22_20_inst : DLH_X1 port map( G => n5148, D => n5022, Q => 
                           registers_22_20_port);
   registers_reg_22_19_inst : DLH_X1 port map( G => n5148, D => n5025, Q => 
                           registers_22_19_port);
   registers_reg_22_18_inst : DLH_X1 port map( G => n5148, D => n5028, Q => 
                           registers_22_18_port);
   registers_reg_22_17_inst : DLH_X1 port map( G => n5148, D => n5031, Q => 
                           registers_22_17_port);
   registers_reg_22_16_inst : DLH_X1 port map( G => n5148, D => n5034, Q => 
                           registers_22_16_port);
   registers_reg_22_15_inst : DLH_X1 port map( G => n5148, D => n5037, Q => 
                           registers_22_15_port);
   registers_reg_22_14_inst : DLH_X1 port map( G => n5148, D => n5040, Q => 
                           registers_22_14_port);
   registers_reg_22_13_inst : DLH_X1 port map( G => n5148, D => n5043, Q => 
                           registers_22_13_port);
   registers_reg_22_12_inst : DLH_X1 port map( G => n5148, D => n5046, Q => 
                           registers_22_12_port);
   registers_reg_22_11_inst : DLH_X1 port map( G => n5148, D => n5049, Q => 
                           registers_22_11_port);
   registers_reg_22_10_inst : DLH_X1 port map( G => n5147, D => n5052, Q => 
                           registers_22_10_port);
   registers_reg_22_9_inst : DLH_X1 port map( G => n5147, D => n5055, Q => 
                           registers_22_9_port);
   registers_reg_22_8_inst : DLH_X1 port map( G => n5147, D => n5058, Q => 
                           registers_22_8_port);
   registers_reg_22_7_inst : DLH_X1 port map( G => n5147, D => n5061, Q => 
                           registers_22_7_port);
   registers_reg_22_6_inst : DLH_X1 port map( G => n5147, D => n5064, Q => 
                           registers_22_6_port);
   registers_reg_22_5_inst : DLH_X1 port map( G => n5147, D => n5067, Q => 
                           registers_22_5_port);
   registers_reg_22_4_inst : DLH_X1 port map( G => n5147, D => n5070, Q => 
                           registers_22_4_port);
   registers_reg_22_3_inst : DLH_X1 port map( G => n5147, D => n5073, Q => 
                           registers_22_3_port);
   registers_reg_22_2_inst : DLH_X1 port map( G => n5147, D => n5076, Q => 
                           registers_22_2_port);
   registers_reg_22_1_inst : DLH_X1 port map( G => n5147, D => n5079, Q => 
                           registers_22_1_port);
   registers_reg_22_0_inst : DLH_X1 port map( G => n5147, D => n5082, Q => 
                           registers_22_0_port);
   registers_reg_23_31_inst : DLH_X1 port map( G => n5152, D => n4988, Q => 
                           registers_23_31_port);
   registers_reg_23_30_inst : DLH_X1 port map( G => n5152, D => n4991, Q => 
                           registers_23_30_port);
   registers_reg_23_29_inst : DLH_X1 port map( G => n5152, D => n4994, Q => 
                           registers_23_29_port);
   registers_reg_23_28_inst : DLH_X1 port map( G => n5152, D => n4997, Q => 
                           registers_23_28_port);
   registers_reg_23_27_inst : DLH_X1 port map( G => n5152, D => n5000, Q => 
                           registers_23_27_port);
   registers_reg_23_26_inst : DLH_X1 port map( G => n5152, D => n5003, Q => 
                           registers_23_26_port);
   registers_reg_23_25_inst : DLH_X1 port map( G => n5152, D => n5006, Q => 
                           registers_23_25_port);
   registers_reg_23_24_inst : DLH_X1 port map( G => n5152, D => n5009, Q => 
                           registers_23_24_port);
   registers_reg_23_23_inst : DLH_X1 port map( G => n5152, D => n5012, Q => 
                           registers_23_23_port);
   registers_reg_23_22_inst : DLH_X1 port map( G => n5152, D => n5015, Q => 
                           registers_23_22_port);
   registers_reg_23_21_inst : DLH_X1 port map( G => n5151, D => n5018, Q => 
                           registers_23_21_port);
   registers_reg_23_20_inst : DLH_X1 port map( G => n5151, D => n5021, Q => 
                           registers_23_20_port);
   registers_reg_23_19_inst : DLH_X1 port map( G => n5151, D => n5024, Q => 
                           registers_23_19_port);
   registers_reg_23_18_inst : DLH_X1 port map( G => n5151, D => n5027, Q => 
                           registers_23_18_port);
   registers_reg_23_17_inst : DLH_X1 port map( G => n5151, D => n5030, Q => 
                           registers_23_17_port);
   registers_reg_23_16_inst : DLH_X1 port map( G => n5151, D => n5033, Q => 
                           registers_23_16_port);
   registers_reg_23_15_inst : DLH_X1 port map( G => n5151, D => n5036, Q => 
                           registers_23_15_port);
   registers_reg_23_14_inst : DLH_X1 port map( G => n5151, D => n5039, Q => 
                           registers_23_14_port);
   registers_reg_23_13_inst : DLH_X1 port map( G => n5151, D => n5042, Q => 
                           registers_23_13_port);
   registers_reg_23_12_inst : DLH_X1 port map( G => n5151, D => n5045, Q => 
                           registers_23_12_port);
   registers_reg_23_11_inst : DLH_X1 port map( G => n5151, D => n5048, Q => 
                           registers_23_11_port);
   registers_reg_23_10_inst : DLH_X1 port map( G => n5150, D => n5051, Q => 
                           registers_23_10_port);
   registers_reg_23_9_inst : DLH_X1 port map( G => n5150, D => n5054, Q => 
                           registers_23_9_port);
   registers_reg_23_8_inst : DLH_X1 port map( G => n5150, D => n5057, Q => 
                           registers_23_8_port);
   registers_reg_23_7_inst : DLH_X1 port map( G => n5150, D => n5060, Q => 
                           registers_23_7_port);
   registers_reg_23_6_inst : DLH_X1 port map( G => n5150, D => n5063, Q => 
                           registers_23_6_port);
   registers_reg_23_5_inst : DLH_X1 port map( G => n5150, D => n5066, Q => 
                           registers_23_5_port);
   registers_reg_23_4_inst : DLH_X1 port map( G => n5150, D => n5069, Q => 
                           registers_23_4_port);
   registers_reg_23_3_inst : DLH_X1 port map( G => n5150, D => n5072, Q => 
                           registers_23_3_port);
   registers_reg_23_2_inst : DLH_X1 port map( G => n5150, D => n5075, Q => 
                           registers_23_2_port);
   registers_reg_23_1_inst : DLH_X1 port map( G => n5150, D => n5078, Q => 
                           registers_23_1_port);
   registers_reg_23_0_inst : DLH_X1 port map( G => n5150, D => n5081, Q => 
                           registers_23_0_port);
   registers_reg_24_31_inst : DLH_X1 port map( G => n5155, D => n4988, Q => 
                           registers_24_31_port);
   registers_reg_24_30_inst : DLH_X1 port map( G => n5155, D => n4991, Q => 
                           registers_24_30_port);
   registers_reg_24_29_inst : DLH_X1 port map( G => n5155, D => n4994, Q => 
                           registers_24_29_port);
   registers_reg_24_28_inst : DLH_X1 port map( G => n5155, D => n4997, Q => 
                           registers_24_28_port);
   registers_reg_24_27_inst : DLH_X1 port map( G => n5155, D => n5000, Q => 
                           registers_24_27_port);
   registers_reg_24_26_inst : DLH_X1 port map( G => n5155, D => n5003, Q => 
                           registers_24_26_port);
   registers_reg_24_25_inst : DLH_X1 port map( G => n5155, D => n5006, Q => 
                           registers_24_25_port);
   registers_reg_24_24_inst : DLH_X1 port map( G => n5155, D => n5009, Q => 
                           registers_24_24_port);
   registers_reg_24_23_inst : DLH_X1 port map( G => n5155, D => n5012, Q => 
                           registers_24_23_port);
   registers_reg_24_22_inst : DLH_X1 port map( G => n5155, D => n5015, Q => 
                           registers_24_22_port);
   registers_reg_24_21_inst : DLH_X1 port map( G => n5154, D => n5018, Q => 
                           registers_24_21_port);
   registers_reg_24_20_inst : DLH_X1 port map( G => n5154, D => n5021, Q => 
                           registers_24_20_port);
   registers_reg_24_19_inst : DLH_X1 port map( G => n5154, D => n5024, Q => 
                           registers_24_19_port);
   registers_reg_24_18_inst : DLH_X1 port map( G => n5154, D => n5027, Q => 
                           registers_24_18_port);
   registers_reg_24_17_inst : DLH_X1 port map( G => n5154, D => n5030, Q => 
                           registers_24_17_port);
   registers_reg_24_16_inst : DLH_X1 port map( G => n5154, D => n5033, Q => 
                           registers_24_16_port);
   registers_reg_24_15_inst : DLH_X1 port map( G => n5154, D => n5036, Q => 
                           registers_24_15_port);
   registers_reg_24_14_inst : DLH_X1 port map( G => n5154, D => n5039, Q => 
                           registers_24_14_port);
   registers_reg_24_13_inst : DLH_X1 port map( G => n5154, D => n5042, Q => 
                           registers_24_13_port);
   registers_reg_24_12_inst : DLH_X1 port map( G => n5154, D => n5045, Q => 
                           registers_24_12_port);
   registers_reg_24_11_inst : DLH_X1 port map( G => n5154, D => n5048, Q => 
                           registers_24_11_port);
   registers_reg_24_10_inst : DLH_X1 port map( G => n5153, D => n5051, Q => 
                           registers_24_10_port);
   registers_reg_24_9_inst : DLH_X1 port map( G => n5153, D => n5054, Q => 
                           registers_24_9_port);
   registers_reg_24_8_inst : DLH_X1 port map( G => n5153, D => n5057, Q => 
                           registers_24_8_port);
   registers_reg_24_7_inst : DLH_X1 port map( G => n5153, D => n5060, Q => 
                           registers_24_7_port);
   registers_reg_24_6_inst : DLH_X1 port map( G => n5153, D => n5063, Q => 
                           registers_24_6_port);
   registers_reg_24_5_inst : DLH_X1 port map( G => n5153, D => n5066, Q => 
                           registers_24_5_port);
   registers_reg_24_4_inst : DLH_X1 port map( G => n5153, D => n5069, Q => 
                           registers_24_4_port);
   registers_reg_24_3_inst : DLH_X1 port map( G => n5153, D => n5072, Q => 
                           registers_24_3_port);
   registers_reg_24_2_inst : DLH_X1 port map( G => n5153, D => n5075, Q => 
                           registers_24_2_port);
   registers_reg_24_1_inst : DLH_X1 port map( G => n5153, D => n5078, Q => 
                           registers_24_1_port);
   registers_reg_24_0_inst : DLH_X1 port map( G => n5153, D => n5081, Q => 
                           registers_24_0_port);
   registers_reg_25_31_inst : DLH_X1 port map( G => n5158, D => n4989, Q => 
                           registers_25_31_port);
   registers_reg_25_30_inst : DLH_X1 port map( G => n5158, D => n4992, Q => 
                           registers_25_30_port);
   registers_reg_25_29_inst : DLH_X1 port map( G => n5158, D => n4995, Q => 
                           registers_25_29_port);
   registers_reg_25_28_inst : DLH_X1 port map( G => n5158, D => n4998, Q => 
                           registers_25_28_port);
   registers_reg_25_27_inst : DLH_X1 port map( G => n5158, D => n5001, Q => 
                           registers_25_27_port);
   registers_reg_25_26_inst : DLH_X1 port map( G => n5158, D => n5004, Q => 
                           registers_25_26_port);
   registers_reg_25_25_inst : DLH_X1 port map( G => n5158, D => n5007, Q => 
                           registers_25_25_port);
   registers_reg_25_24_inst : DLH_X1 port map( G => n5158, D => n5010, Q => 
                           registers_25_24_port);
   registers_reg_25_23_inst : DLH_X1 port map( G => n5158, D => n5013, Q => 
                           registers_25_23_port);
   registers_reg_25_22_inst : DLH_X1 port map( G => n5158, D => n5016, Q => 
                           registers_25_22_port);
   registers_reg_25_21_inst : DLH_X1 port map( G => n5157, D => n5019, Q => 
                           registers_25_21_port);
   registers_reg_25_20_inst : DLH_X1 port map( G => n5157, D => n5022, Q => 
                           registers_25_20_port);
   registers_reg_25_19_inst : DLH_X1 port map( G => n5157, D => n5025, Q => 
                           registers_25_19_port);
   registers_reg_25_18_inst : DLH_X1 port map( G => n5157, D => n5028, Q => 
                           registers_25_18_port);
   registers_reg_25_17_inst : DLH_X1 port map( G => n5157, D => n5031, Q => 
                           registers_25_17_port);
   registers_reg_25_16_inst : DLH_X1 port map( G => n5157, D => n5034, Q => 
                           registers_25_16_port);
   registers_reg_25_15_inst : DLH_X1 port map( G => n5157, D => n5037, Q => 
                           registers_25_15_port);
   registers_reg_25_14_inst : DLH_X1 port map( G => n5157, D => n5040, Q => 
                           registers_25_14_port);
   registers_reg_25_13_inst : DLH_X1 port map( G => n5157, D => n5043, Q => 
                           registers_25_13_port);
   registers_reg_25_12_inst : DLH_X1 port map( G => n5157, D => n5046, Q => 
                           registers_25_12_port);
   registers_reg_25_11_inst : DLH_X1 port map( G => n5157, D => n5049, Q => 
                           registers_25_11_port);
   registers_reg_25_10_inst : DLH_X1 port map( G => n5156, D => n5052, Q => 
                           registers_25_10_port);
   registers_reg_25_9_inst : DLH_X1 port map( G => n5156, D => n5055, Q => 
                           registers_25_9_port);
   registers_reg_25_8_inst : DLH_X1 port map( G => n5156, D => n5058, Q => 
                           registers_25_8_port);
   registers_reg_25_7_inst : DLH_X1 port map( G => n5156, D => n5061, Q => 
                           registers_25_7_port);
   registers_reg_25_6_inst : DLH_X1 port map( G => n5156, D => n5064, Q => 
                           registers_25_6_port);
   registers_reg_25_5_inst : DLH_X1 port map( G => n5156, D => n5067, Q => 
                           registers_25_5_port);
   registers_reg_25_4_inst : DLH_X1 port map( G => n5156, D => n5070, Q => 
                           registers_25_4_port);
   registers_reg_25_3_inst : DLH_X1 port map( G => n5156, D => n5073, Q => 
                           registers_25_3_port);
   registers_reg_25_2_inst : DLH_X1 port map( G => n5156, D => n5076, Q => 
                           registers_25_2_port);
   registers_reg_25_1_inst : DLH_X1 port map( G => n5156, D => n5079, Q => 
                           registers_25_1_port);
   registers_reg_25_0_inst : DLH_X1 port map( G => n5156, D => n5082, Q => 
                           registers_25_0_port);
   registers_reg_26_31_inst : DLH_X1 port map( G => n5161, D => n4989, Q => 
                           registers_26_31_port);
   registers_reg_26_30_inst : DLH_X1 port map( G => n5161, D => n4992, Q => 
                           registers_26_30_port);
   registers_reg_26_29_inst : DLH_X1 port map( G => n5161, D => n4995, Q => 
                           registers_26_29_port);
   registers_reg_26_28_inst : DLH_X1 port map( G => n5161, D => n4998, Q => 
                           registers_26_28_port);
   registers_reg_26_27_inst : DLH_X1 port map( G => n5161, D => n5001, Q => 
                           registers_26_27_port);
   registers_reg_26_26_inst : DLH_X1 port map( G => n5161, D => n5004, Q => 
                           registers_26_26_port);
   registers_reg_26_25_inst : DLH_X1 port map( G => n5161, D => n5007, Q => 
                           registers_26_25_port);
   registers_reg_26_24_inst : DLH_X1 port map( G => n5161, D => n5010, Q => 
                           registers_26_24_port);
   registers_reg_26_23_inst : DLH_X1 port map( G => n5161, D => n5013, Q => 
                           registers_26_23_port);
   registers_reg_26_22_inst : DLH_X1 port map( G => n5161, D => n5016, Q => 
                           registers_26_22_port);
   registers_reg_26_21_inst : DLH_X1 port map( G => n5160, D => n5019, Q => 
                           registers_26_21_port);
   registers_reg_26_20_inst : DLH_X1 port map( G => n5160, D => n5022, Q => 
                           registers_26_20_port);
   registers_reg_26_19_inst : DLH_X1 port map( G => n5160, D => n5025, Q => 
                           registers_26_19_port);
   registers_reg_26_18_inst : DLH_X1 port map( G => n5160, D => n5028, Q => 
                           registers_26_18_port);
   registers_reg_26_17_inst : DLH_X1 port map( G => n5160, D => n5031, Q => 
                           registers_26_17_port);
   registers_reg_26_16_inst : DLH_X1 port map( G => n5160, D => n5034, Q => 
                           registers_26_16_port);
   registers_reg_26_15_inst : DLH_X1 port map( G => n5160, D => n5037, Q => 
                           registers_26_15_port);
   registers_reg_26_14_inst : DLH_X1 port map( G => n5160, D => n5040, Q => 
                           registers_26_14_port);
   registers_reg_26_13_inst : DLH_X1 port map( G => n5160, D => n5043, Q => 
                           registers_26_13_port);
   registers_reg_26_12_inst : DLH_X1 port map( G => n5160, D => n5046, Q => 
                           registers_26_12_port);
   registers_reg_26_11_inst : DLH_X1 port map( G => n5160, D => n5049, Q => 
                           registers_26_11_port);
   registers_reg_26_10_inst : DLH_X1 port map( G => n5159, D => n5052, Q => 
                           registers_26_10_port);
   registers_reg_26_9_inst : DLH_X1 port map( G => n5159, D => n5055, Q => 
                           registers_26_9_port);
   registers_reg_26_8_inst : DLH_X1 port map( G => n5159, D => n5058, Q => 
                           registers_26_8_port);
   registers_reg_26_7_inst : DLH_X1 port map( G => n5159, D => n5061, Q => 
                           registers_26_7_port);
   registers_reg_26_6_inst : DLH_X1 port map( G => n5159, D => n5064, Q => 
                           registers_26_6_port);
   registers_reg_26_5_inst : DLH_X1 port map( G => n5159, D => n5067, Q => 
                           registers_26_5_port);
   registers_reg_26_4_inst : DLH_X1 port map( G => n5159, D => n5070, Q => 
                           registers_26_4_port);
   registers_reg_26_3_inst : DLH_X1 port map( G => n5159, D => n5073, Q => 
                           registers_26_3_port);
   registers_reg_26_2_inst : DLH_X1 port map( G => n5159, D => n5076, Q => 
                           registers_26_2_port);
   registers_reg_26_1_inst : DLH_X1 port map( G => n5159, D => n5079, Q => 
                           registers_26_1_port);
   registers_reg_26_0_inst : DLH_X1 port map( G => n5159, D => n5082, Q => 
                           registers_26_0_port);
   registers_reg_27_31_inst : DLH_X1 port map( G => n5164, D => n4989, Q => 
                           registers_27_31_port);
   registers_reg_27_30_inst : DLH_X1 port map( G => n5164, D => n4992, Q => 
                           registers_27_30_port);
   registers_reg_27_29_inst : DLH_X1 port map( G => n5164, D => n4995, Q => 
                           registers_27_29_port);
   registers_reg_27_28_inst : DLH_X1 port map( G => n5164, D => n4998, Q => 
                           registers_27_28_port);
   registers_reg_27_27_inst : DLH_X1 port map( G => n5164, D => n5001, Q => 
                           registers_27_27_port);
   registers_reg_27_26_inst : DLH_X1 port map( G => n5164, D => n5004, Q => 
                           registers_27_26_port);
   registers_reg_27_25_inst : DLH_X1 port map( G => n5164, D => n5007, Q => 
                           registers_27_25_port);
   registers_reg_27_24_inst : DLH_X1 port map( G => n5164, D => n5010, Q => 
                           registers_27_24_port);
   registers_reg_27_23_inst : DLH_X1 port map( G => n5164, D => n5013, Q => 
                           registers_27_23_port);
   registers_reg_27_22_inst : DLH_X1 port map( G => n5164, D => n5016, Q => 
                           registers_27_22_port);
   registers_reg_27_21_inst : DLH_X1 port map( G => n5163, D => n5019, Q => 
                           registers_27_21_port);
   registers_reg_27_20_inst : DLH_X1 port map( G => n5163, D => n5022, Q => 
                           registers_27_20_port);
   registers_reg_27_19_inst : DLH_X1 port map( G => n5163, D => n5025, Q => 
                           registers_27_19_port);
   registers_reg_27_18_inst : DLH_X1 port map( G => n5163, D => n5028, Q => 
                           registers_27_18_port);
   registers_reg_27_17_inst : DLH_X1 port map( G => n5163, D => n5031, Q => 
                           registers_27_17_port);
   registers_reg_27_16_inst : DLH_X1 port map( G => n5163, D => n5034, Q => 
                           registers_27_16_port);
   registers_reg_27_15_inst : DLH_X1 port map( G => n5163, D => n5037, Q => 
                           registers_27_15_port);
   registers_reg_27_14_inst : DLH_X1 port map( G => n5163, D => n5040, Q => 
                           registers_27_14_port);
   registers_reg_27_13_inst : DLH_X1 port map( G => n5163, D => n5043, Q => 
                           registers_27_13_port);
   registers_reg_27_12_inst : DLH_X1 port map( G => n5163, D => n5046, Q => 
                           registers_27_12_port);
   registers_reg_27_11_inst : DLH_X1 port map( G => n5163, D => n5049, Q => 
                           registers_27_11_port);
   registers_reg_27_10_inst : DLH_X1 port map( G => n5162, D => n5052, Q => 
                           registers_27_10_port);
   registers_reg_27_9_inst : DLH_X1 port map( G => n5162, D => n5055, Q => 
                           registers_27_9_port);
   registers_reg_27_8_inst : DLH_X1 port map( G => n5162, D => n5058, Q => 
                           registers_27_8_port);
   registers_reg_27_7_inst : DLH_X1 port map( G => n5162, D => n5061, Q => 
                           registers_27_7_port);
   registers_reg_27_6_inst : DLH_X1 port map( G => n5162, D => n5064, Q => 
                           registers_27_6_port);
   registers_reg_27_5_inst : DLH_X1 port map( G => n5162, D => n5067, Q => 
                           registers_27_5_port);
   registers_reg_27_4_inst : DLH_X1 port map( G => n5162, D => n5070, Q => 
                           registers_27_4_port);
   registers_reg_27_3_inst : DLH_X1 port map( G => n5162, D => n5073, Q => 
                           registers_27_3_port);
   registers_reg_27_2_inst : DLH_X1 port map( G => n5162, D => n5076, Q => 
                           registers_27_2_port);
   registers_reg_27_1_inst : DLH_X1 port map( G => n5162, D => n5079, Q => 
                           registers_27_1_port);
   registers_reg_27_0_inst : DLH_X1 port map( G => n5162, D => n5082, Q => 
                           registers_27_0_port);
   registers_reg_28_31_inst : DLH_X1 port map( G => n5167, D => n4989, Q => 
                           registers_28_31_port);
   registers_reg_28_30_inst : DLH_X1 port map( G => n5167, D => n4992, Q => 
                           registers_28_30_port);
   registers_reg_28_29_inst : DLH_X1 port map( G => n5167, D => n4995, Q => 
                           registers_28_29_port);
   registers_reg_28_28_inst : DLH_X1 port map( G => n5167, D => n4998, Q => 
                           registers_28_28_port);
   registers_reg_28_27_inst : DLH_X1 port map( G => n5167, D => n5001, Q => 
                           registers_28_27_port);
   registers_reg_28_26_inst : DLH_X1 port map( G => n5167, D => n5004, Q => 
                           registers_28_26_port);
   registers_reg_28_25_inst : DLH_X1 port map( G => n5167, D => n5007, Q => 
                           registers_28_25_port);
   registers_reg_28_24_inst : DLH_X1 port map( G => n5167, D => n5010, Q => 
                           registers_28_24_port);
   registers_reg_28_23_inst : DLH_X1 port map( G => n5167, D => n5013, Q => 
                           registers_28_23_port);
   registers_reg_28_22_inst : DLH_X1 port map( G => n5167, D => n5016, Q => 
                           registers_28_22_port);
   registers_reg_28_21_inst : DLH_X1 port map( G => n5166, D => n5019, Q => 
                           registers_28_21_port);
   registers_reg_28_20_inst : DLH_X1 port map( G => n5166, D => n5022, Q => 
                           registers_28_20_port);
   registers_reg_28_19_inst : DLH_X1 port map( G => n5166, D => n5025, Q => 
                           registers_28_19_port);
   registers_reg_28_18_inst : DLH_X1 port map( G => n5166, D => n5028, Q => 
                           registers_28_18_port);
   registers_reg_28_17_inst : DLH_X1 port map( G => n5166, D => n5031, Q => 
                           registers_28_17_port);
   registers_reg_28_16_inst : DLH_X1 port map( G => n5166, D => n5034, Q => 
                           registers_28_16_port);
   registers_reg_28_15_inst : DLH_X1 port map( G => n5166, D => n5037, Q => 
                           registers_28_15_port);
   registers_reg_28_14_inst : DLH_X1 port map( G => n5166, D => n5040, Q => 
                           registers_28_14_port);
   registers_reg_28_13_inst : DLH_X1 port map( G => n5166, D => n5043, Q => 
                           registers_28_13_port);
   registers_reg_28_12_inst : DLH_X1 port map( G => n5166, D => n5046, Q => 
                           registers_28_12_port);
   registers_reg_28_11_inst : DLH_X1 port map( G => n5166, D => n5049, Q => 
                           registers_28_11_port);
   registers_reg_28_10_inst : DLH_X1 port map( G => n5165, D => n5052, Q => 
                           registers_28_10_port);
   registers_reg_28_9_inst : DLH_X1 port map( G => n5165, D => n5055, Q => 
                           registers_28_9_port);
   registers_reg_28_8_inst : DLH_X1 port map( G => n5165, D => n5058, Q => 
                           registers_28_8_port);
   registers_reg_28_7_inst : DLH_X1 port map( G => n5165, D => n5061, Q => 
                           registers_28_7_port);
   registers_reg_28_6_inst : DLH_X1 port map( G => n5165, D => n5064, Q => 
                           registers_28_6_port);
   registers_reg_28_5_inst : DLH_X1 port map( G => n5165, D => n5067, Q => 
                           registers_28_5_port);
   registers_reg_28_4_inst : DLH_X1 port map( G => n5165, D => n5070, Q => 
                           registers_28_4_port);
   registers_reg_28_3_inst : DLH_X1 port map( G => n5165, D => n5073, Q => 
                           registers_28_3_port);
   registers_reg_28_2_inst : DLH_X1 port map( G => n5165, D => n5076, Q => 
                           registers_28_2_port);
   registers_reg_28_1_inst : DLH_X1 port map( G => n5165, D => n5079, Q => 
                           registers_28_1_port);
   registers_reg_28_0_inst : DLH_X1 port map( G => n5165, D => n5082, Q => 
                           registers_28_0_port);
   registers_reg_29_31_inst : DLH_X1 port map( G => n5170, D => n4989, Q => 
                           registers_29_31_port);
   registers_reg_29_30_inst : DLH_X1 port map( G => n5170, D => n4992, Q => 
                           registers_29_30_port);
   registers_reg_29_29_inst : DLH_X1 port map( G => n5170, D => n4995, Q => 
                           registers_29_29_port);
   registers_reg_29_28_inst : DLH_X1 port map( G => n5170, D => n4998, Q => 
                           registers_29_28_port);
   registers_reg_29_27_inst : DLH_X1 port map( G => n5170, D => n5001, Q => 
                           registers_29_27_port);
   registers_reg_29_26_inst : DLH_X1 port map( G => n5170, D => n5004, Q => 
                           registers_29_26_port);
   registers_reg_29_25_inst : DLH_X1 port map( G => n5170, D => n5007, Q => 
                           registers_29_25_port);
   registers_reg_29_24_inst : DLH_X1 port map( G => n5170, D => n5010, Q => 
                           registers_29_24_port);
   registers_reg_29_23_inst : DLH_X1 port map( G => n5170, D => n5013, Q => 
                           registers_29_23_port);
   registers_reg_29_22_inst : DLH_X1 port map( G => n5170, D => n5016, Q => 
                           registers_29_22_port);
   registers_reg_29_21_inst : DLH_X1 port map( G => n5169, D => n5019, Q => 
                           registers_29_21_port);
   registers_reg_29_20_inst : DLH_X1 port map( G => n5169, D => n5022, Q => 
                           registers_29_20_port);
   registers_reg_29_19_inst : DLH_X1 port map( G => n5169, D => n5025, Q => 
                           registers_29_19_port);
   registers_reg_29_18_inst : DLH_X1 port map( G => n5169, D => n5028, Q => 
                           registers_29_18_port);
   registers_reg_29_17_inst : DLH_X1 port map( G => n5169, D => n5031, Q => 
                           registers_29_17_port);
   registers_reg_29_16_inst : DLH_X1 port map( G => n5169, D => n5034, Q => 
                           registers_29_16_port);
   registers_reg_29_15_inst : DLH_X1 port map( G => n5169, D => n5037, Q => 
                           registers_29_15_port);
   registers_reg_29_14_inst : DLH_X1 port map( G => n5169, D => n5040, Q => 
                           registers_29_14_port);
   registers_reg_29_13_inst : DLH_X1 port map( G => n5169, D => n5043, Q => 
                           registers_29_13_port);
   registers_reg_29_12_inst : DLH_X1 port map( G => n5169, D => n5046, Q => 
                           registers_29_12_port);
   registers_reg_29_11_inst : DLH_X1 port map( G => n5169, D => n5049, Q => 
                           registers_29_11_port);
   registers_reg_29_10_inst : DLH_X1 port map( G => n5168, D => n5052, Q => 
                           registers_29_10_port);
   registers_reg_29_9_inst : DLH_X1 port map( G => n5168, D => n5055, Q => 
                           registers_29_9_port);
   registers_reg_29_8_inst : DLH_X1 port map( G => n5168, D => n5058, Q => 
                           registers_29_8_port);
   registers_reg_29_7_inst : DLH_X1 port map( G => n5168, D => n5061, Q => 
                           registers_29_7_port);
   registers_reg_29_6_inst : DLH_X1 port map( G => n5168, D => n5064, Q => 
                           registers_29_6_port);
   registers_reg_29_5_inst : DLH_X1 port map( G => n5168, D => n5067, Q => 
                           registers_29_5_port);
   registers_reg_29_4_inst : DLH_X1 port map( G => n5168, D => n5070, Q => 
                           registers_29_4_port);
   registers_reg_29_3_inst : DLH_X1 port map( G => n5168, D => n5073, Q => 
                           registers_29_3_port);
   registers_reg_29_2_inst : DLH_X1 port map( G => n5168, D => n5076, Q => 
                           registers_29_2_port);
   registers_reg_29_1_inst : DLH_X1 port map( G => n5168, D => n5079, Q => 
                           registers_29_1_port);
   registers_reg_29_0_inst : DLH_X1 port map( G => n5168, D => n5082, Q => 
                           registers_29_0_port);
   registers_reg_30_31_inst : DLH_X1 port map( G => n5173, D => n4989, Q => 
                           registers_30_31_port);
   registers_reg_30_30_inst : DLH_X1 port map( G => n5173, D => n4992, Q => 
                           registers_30_30_port);
   registers_reg_30_29_inst : DLH_X1 port map( G => n5173, D => n4995, Q => 
                           registers_30_29_port);
   registers_reg_30_28_inst : DLH_X1 port map( G => n5173, D => n4998, Q => 
                           registers_30_28_port);
   registers_reg_30_27_inst : DLH_X1 port map( G => n5173, D => n5001, Q => 
                           registers_30_27_port);
   registers_reg_30_26_inst : DLH_X1 port map( G => n5173, D => n5004, Q => 
                           registers_30_26_port);
   registers_reg_30_25_inst : DLH_X1 port map( G => n5173, D => n5007, Q => 
                           registers_30_25_port);
   registers_reg_30_24_inst : DLH_X1 port map( G => n5173, D => n5010, Q => 
                           registers_30_24_port);
   registers_reg_30_23_inst : DLH_X1 port map( G => n5173, D => n5013, Q => 
                           registers_30_23_port);
   registers_reg_30_22_inst : DLH_X1 port map( G => n5173, D => n5016, Q => 
                           registers_30_22_port);
   registers_reg_30_21_inst : DLH_X1 port map( G => n5172, D => n5019, Q => 
                           registers_30_21_port);
   registers_reg_30_20_inst : DLH_X1 port map( G => n5172, D => n5022, Q => 
                           registers_30_20_port);
   registers_reg_30_19_inst : DLH_X1 port map( G => n5172, D => n5025, Q => 
                           registers_30_19_port);
   registers_reg_30_18_inst : DLH_X1 port map( G => n5172, D => n5028, Q => 
                           registers_30_18_port);
   registers_reg_30_17_inst : DLH_X1 port map( G => n5172, D => n5031, Q => 
                           registers_30_17_port);
   registers_reg_30_16_inst : DLH_X1 port map( G => n5172, D => n5034, Q => 
                           registers_30_16_port);
   registers_reg_30_15_inst : DLH_X1 port map( G => n5172, D => n5037, Q => 
                           registers_30_15_port);
   registers_reg_30_14_inst : DLH_X1 port map( G => n5172, D => n5040, Q => 
                           registers_30_14_port);
   registers_reg_30_13_inst : DLH_X1 port map( G => n5172, D => n5043, Q => 
                           registers_30_13_port);
   registers_reg_30_12_inst : DLH_X1 port map( G => n5172, D => n5046, Q => 
                           registers_30_12_port);
   registers_reg_30_11_inst : DLH_X1 port map( G => n5172, D => n5049, Q => 
                           registers_30_11_port);
   registers_reg_30_10_inst : DLH_X1 port map( G => n5171, D => n5052, Q => 
                           registers_30_10_port);
   registers_reg_30_9_inst : DLH_X1 port map( G => n5171, D => n5055, Q => 
                           registers_30_9_port);
   registers_reg_30_8_inst : DLH_X1 port map( G => n5171, D => n5058, Q => 
                           registers_30_8_port);
   registers_reg_30_7_inst : DLH_X1 port map( G => n5171, D => n5061, Q => 
                           registers_30_7_port);
   registers_reg_30_6_inst : DLH_X1 port map( G => n5171, D => n5064, Q => 
                           registers_30_6_port);
   registers_reg_30_5_inst : DLH_X1 port map( G => n5171, D => n5067, Q => 
                           registers_30_5_port);
   registers_reg_30_4_inst : DLH_X1 port map( G => n5171, D => n5070, Q => 
                           registers_30_4_port);
   registers_reg_30_3_inst : DLH_X1 port map( G => n5171, D => n5073, Q => 
                           registers_30_3_port);
   registers_reg_30_2_inst : DLH_X1 port map( G => n5171, D => n5076, Q => 
                           registers_30_2_port);
   registers_reg_30_1_inst : DLH_X1 port map( G => n5171, D => n5079, Q => 
                           registers_30_1_port);
   registers_reg_30_0_inst : DLH_X1 port map( G => n5171, D => n5082, Q => 
                           registers_30_0_port);
   registers_reg_31_31_inst : DLH_X1 port map( G => n5176, D => n4989, Q => 
                           registers_31_31_port);
   registers_reg_31_30_inst : DLH_X1 port map( G => n5176, D => n4992, Q => 
                           registers_31_30_port);
   registers_reg_31_29_inst : DLH_X1 port map( G => n5176, D => n4995, Q => 
                           registers_31_29_port);
   registers_reg_31_28_inst : DLH_X1 port map( G => n5176, D => n4998, Q => 
                           registers_31_28_port);
   registers_reg_31_27_inst : DLH_X1 port map( G => n5176, D => n5001, Q => 
                           registers_31_27_port);
   registers_reg_31_26_inst : DLH_X1 port map( G => n5176, D => n5004, Q => 
                           registers_31_26_port);
   registers_reg_31_25_inst : DLH_X1 port map( G => n5176, D => n5007, Q => 
                           registers_31_25_port);
   registers_reg_31_24_inst : DLH_X1 port map( G => n5176, D => n5010, Q => 
                           registers_31_24_port);
   registers_reg_31_23_inst : DLH_X1 port map( G => n5176, D => n5013, Q => 
                           registers_31_23_port);
   registers_reg_31_22_inst : DLH_X1 port map( G => n5176, D => n5016, Q => 
                           registers_31_22_port);
   registers_reg_31_21_inst : DLH_X1 port map( G => n5175, D => n5019, Q => 
                           registers_31_21_port);
   registers_reg_31_20_inst : DLH_X1 port map( G => n5175, D => n5022, Q => 
                           registers_31_20_port);
   registers_reg_31_19_inst : DLH_X1 port map( G => n5175, D => n5025, Q => 
                           registers_31_19_port);
   registers_reg_31_18_inst : DLH_X1 port map( G => n5175, D => n5028, Q => 
                           registers_31_18_port);
   registers_reg_31_17_inst : DLH_X1 port map( G => n5175, D => n5031, Q => 
                           registers_31_17_port);
   registers_reg_31_16_inst : DLH_X1 port map( G => n5175, D => n5034, Q => 
                           registers_31_16_port);
   registers_reg_31_15_inst : DLH_X1 port map( G => n5175, D => n5037, Q => 
                           registers_31_15_port);
   registers_reg_31_14_inst : DLH_X1 port map( G => n5175, D => n5040, Q => 
                           registers_31_14_port);
   registers_reg_31_13_inst : DLH_X1 port map( G => n5175, D => n5043, Q => 
                           registers_31_13_port);
   registers_reg_31_12_inst : DLH_X1 port map( G => n5175, D => n5046, Q => 
                           registers_31_12_port);
   registers_reg_31_11_inst : DLH_X1 port map( G => n5175, D => n5049, Q => 
                           registers_31_11_port);
   registers_reg_31_10_inst : DLH_X1 port map( G => n5174, D => n5052, Q => 
                           registers_31_10_port);
   registers_reg_31_9_inst : DLH_X1 port map( G => n5174, D => n5055, Q => 
                           registers_31_9_port);
   registers_reg_31_8_inst : DLH_X1 port map( G => n5174, D => n5058, Q => 
                           registers_31_8_port);
   registers_reg_31_7_inst : DLH_X1 port map( G => n5174, D => n5061, Q => 
                           registers_31_7_port);
   registers_reg_31_6_inst : DLH_X1 port map( G => n5174, D => n5064, Q => 
                           registers_31_6_port);
   registers_reg_31_5_inst : DLH_X1 port map( G => n5174, D => n5067, Q => 
                           registers_31_5_port);
   registers_reg_31_4_inst : DLH_X1 port map( G => n5174, D => n5070, Q => 
                           registers_31_4_port);
   registers_reg_31_3_inst : DLH_X1 port map( G => n5174, D => n5073, Q => 
                           registers_31_3_port);
   registers_reg_31_2_inst : DLH_X1 port map( G => n5174, D => n5076, Q => 
                           registers_31_2_port);
   registers_reg_31_1_inst : DLH_X1 port map( G => n5174, D => n5079, Q => 
                           registers_31_1_port);
   registers_reg_31_0_inst : DLH_X1 port map( G => n5174, D => n5082, Q => 
                           registers_31_0_port);
   U1834 : NAND3_X1 port map( A1 => n538, A2 => n539, A3 => w_signal, ZN => 
                           n530);
   U1835 : NAND3_X1 port map( A1 => w_signal, A2 => n539, A3 => 
                           address_port_w(3), ZN => n540);
   U1836 : NAND3_X1 port map( A1 => w_signal, A2 => n538, A3 => 
                           address_port_w(4), ZN => n542);
   U1837 : NAND3_X1 port map( A1 => n544, A2 => n545, A3 => n546, ZN => n541);
   U1838 : NAND3_X1 port map( A1 => n544, A2 => n545, A3 => address_port_w(0), 
                           ZN => n531);
   U1839 : NAND3_X1 port map( A1 => n546, A2 => n545, A3 => address_port_w(1), 
                           ZN => n532);
   U1840 : NAND3_X1 port map( A1 => address_port_w(0), A2 => n545, A3 => 
                           address_port_w(1), ZN => n533);
   U1841 : NAND3_X1 port map( A1 => n546, A2 => n544, A3 => address_port_w(2), 
                           ZN => n534);
   U1842 : NAND3_X1 port map( A1 => address_port_w(0), A2 => n544, A3 => 
                           address_port_w(2), ZN => n535);
   U1843 : NAND3_X1 port map( A1 => address_port_w(1), A2 => n546, A3 => 
                           address_port_w(2), ZN => n536);
   U1844 : NAND3_X1 port map( A1 => address_port_w(3), A2 => w_signal, A3 => 
                           address_port_w(4), ZN => n543);
   U1845 : NAND3_X1 port map( A1 => address_port_w(1), A2 => address_port_w(0),
                           A3 => address_port_w(2), ZN => n537);
   data_out_port_a_tri_24_inst : TBUF_X1 port map( A => n1818, EN => n4983, Z 
                           => data_out_port_a(24));
   data_out_port_a_tri_25_inst : TBUF_X1 port map( A => n1817, EN => n4983, Z 
                           => data_out_port_a(25));
   data_out_port_a_tri_26_inst : TBUF_X1 port map( A => n1816, EN => n4983, Z 
                           => data_out_port_a(26));
   data_out_port_a_tri_27_inst : TBUF_X1 port map( A => n1815, EN => n4983, Z 
                           => data_out_port_a(27));
   data_out_port_a_tri_28_inst : TBUF_X1 port map( A => n1814, EN => n4983, Z 
                           => data_out_port_a(28));
   data_out_port_a_tri_29_inst : TBUF_X1 port map( A => n1813, EN => n4983, Z 
                           => data_out_port_a(29));
   data_out_port_a_tri_30_inst : TBUF_X1 port map( A => n1812, EN => n4983, Z 
                           => data_out_port_a(30));
   data_out_port_a_tri_31_inst : TBUF_X1 port map( A => n1811, EN => n4983, Z 
                           => data_out_port_a(31));
   data_out_port_b_tri_24_inst : TBUF_X1 port map( A => n1785, EN => n4986, Z 
                           => data_out_port_b(24));
   data_out_port_b_tri_25_inst : TBUF_X1 port map( A => n1784, EN => n4986, Z 
                           => data_out_port_b(25));
   data_out_port_b_tri_26_inst : TBUF_X1 port map( A => n1783, EN => n4986, Z 
                           => data_out_port_b(26));
   data_out_port_b_tri_27_inst : TBUF_X1 port map( A => n1782, EN => n4986, Z 
                           => data_out_port_b(27));
   data_out_port_b_tri_28_inst : TBUF_X1 port map( A => n1781, EN => n4986, Z 
                           => data_out_port_b(28));
   data_out_port_b_tri_29_inst : TBUF_X1 port map( A => n1780, EN => n4986, Z 
                           => data_out_port_b(29));
   data_out_port_b_tri_30_inst : TBUF_X1 port map( A => n1779, EN => n4986, Z 
                           => data_out_port_b(30));
   data_out_port_b_tri_31_inst : TBUF_X1 port map( A => n1778, EN => n4986, Z 
                           => data_out_port_b(31));
   data_out_port_a_tri_0_inst : TBUF_X1 port map( A => n1843, EN => n4983, Z =>
                           data_out_port_a(0));
   data_out_port_a_tri_1_inst : TBUF_X1 port map( A => n1842, EN => n4983, Z =>
                           data_out_port_a(1));
   data_out_port_a_tri_2_inst : TBUF_X1 port map( A => n1841, EN => n4983, Z =>
                           data_out_port_a(2));
   data_out_port_a_tri_3_inst : TBUF_X1 port map( A => n1840, EN => n4983, Z =>
                           data_out_port_a(3));
   data_out_port_a_tri_4_inst : TBUF_X1 port map( A => n1839, EN => n4982, Z =>
                           data_out_port_a(4));
   data_out_port_a_tri_5_inst : TBUF_X1 port map( A => n1838, EN => n4982, Z =>
                           data_out_port_a(5));
   data_out_port_a_tri_6_inst : TBUF_X1 port map( A => n1837, EN => n4982, Z =>
                           data_out_port_a(6));
   data_out_port_a_tri_7_inst : TBUF_X1 port map( A => n1836, EN => n4982, Z =>
                           data_out_port_a(7));
   data_out_port_b_tri_0_inst : TBUF_X1 port map( A => n1810, EN => n4986, Z =>
                           data_out_port_b(0));
   data_out_port_b_tri_1_inst : TBUF_X1 port map( A => n1809, EN => n4986, Z =>
                           data_out_port_b(1));
   data_out_port_b_tri_2_inst : TBUF_X1 port map( A => n1808, EN => n4986, Z =>
                           data_out_port_b(2));
   data_out_port_b_tri_3_inst : TBUF_X1 port map( A => n1807, EN => n4986, Z =>
                           data_out_port_b(3));
   data_out_port_b_tri_4_inst : TBUF_X1 port map( A => n1806, EN => n4985, Z =>
                           data_out_port_b(4));
   data_out_port_b_tri_5_inst : TBUF_X1 port map( A => n1805, EN => n4985, Z =>
                           data_out_port_b(5));
   data_out_port_b_tri_6_inst : TBUF_X1 port map( A => n1804, EN => n4985, Z =>
                           data_out_port_b(6));
   data_out_port_b_tri_7_inst : TBUF_X1 port map( A => n1803, EN => n4985, Z =>
                           data_out_port_b(7));
   data_out_port_a_tri_8_inst : TBUF_X1 port map( A => n1835, EN => n4982, Z =>
                           data_out_port_a(8));
   data_out_port_a_tri_9_inst : TBUF_X1 port map( A => n1833, EN => n4982, Z =>
                           data_out_port_a(9));
   data_out_port_a_tri_10_inst : TBUF_X1 port map( A => n1832, EN => n4982, Z 
                           => data_out_port_a(10));
   data_out_port_a_tri_11_inst : TBUF_X1 port map( A => n1831, EN => n4982, Z 
                           => data_out_port_a(11));
   data_out_port_a_tri_12_inst : TBUF_X1 port map( A => n1830, EN => n4982, Z 
                           => data_out_port_a(12));
   data_out_port_a_tri_13_inst : TBUF_X1 port map( A => n1829, EN => n4982, Z 
                           => data_out_port_a(13));
   data_out_port_a_tri_14_inst : TBUF_X1 port map( A => n1828, EN => n4982, Z 
                           => data_out_port_a(14));
   data_out_port_a_tri_15_inst : TBUF_X1 port map( A => n1827, EN => n4982, Z 
                           => data_out_port_a(15));
   data_out_port_b_tri_8_inst : TBUF_X1 port map( A => n1802, EN => n4985, Z =>
                           data_out_port_b(8));
   data_out_port_b_tri_9_inst : TBUF_X1 port map( A => n1800, EN => n4985, Z =>
                           data_out_port_b(9));
   data_out_port_b_tri_10_inst : TBUF_X1 port map( A => n1799, EN => n4985, Z 
                           => data_out_port_b(10));
   data_out_port_b_tri_11_inst : TBUF_X1 port map( A => n1798, EN => n4985, Z 
                           => data_out_port_b(11));
   data_out_port_b_tri_12_inst : TBUF_X1 port map( A => n1797, EN => n4985, Z 
                           => data_out_port_b(12));
   data_out_port_b_tri_13_inst : TBUF_X1 port map( A => n1796, EN => n4985, Z 
                           => data_out_port_b(13));
   data_out_port_b_tri_14_inst : TBUF_X1 port map( A => n1795, EN => n4985, Z 
                           => data_out_port_b(14));
   data_out_port_b_tri_15_inst : TBUF_X1 port map( A => n1794, EN => n4985, Z 
                           => data_out_port_b(15));
   data_out_port_a_tri_16_inst : TBUF_X1 port map( A => n1826, EN => n4984, Z 
                           => data_out_port_a(16));
   data_out_port_a_tri_17_inst : TBUF_X1 port map( A => n1825, EN => n4984, Z 
                           => data_out_port_a(17));
   data_out_port_a_tri_18_inst : TBUF_X1 port map( A => n1824, EN => n4984, Z 
                           => data_out_port_a(18));
   data_out_port_a_tri_19_inst : TBUF_X1 port map( A => n1823, EN => n4984, Z 
                           => data_out_port_a(19));
   data_out_port_a_tri_20_inst : TBUF_X1 port map( A => n1822, EN => n4984, Z 
                           => data_out_port_a(20));
   data_out_port_a_tri_21_inst : TBUF_X1 port map( A => n1821, EN => n4984, Z 
                           => data_out_port_a(21));
   data_out_port_a_tri_22_inst : TBUF_X1 port map( A => n1820, EN => n4984, Z 
                           => data_out_port_a(22));
   data_out_port_a_tri_23_inst : TBUF_X1 port map( A => n1819, EN => n4984, Z 
                           => data_out_port_a(23));
   data_out_port_b_tri_16_inst : TBUF_X1 port map( A => n1793, EN => n4987, Z 
                           => data_out_port_b(16));
   data_out_port_b_tri_17_inst : TBUF_X1 port map( A => n1792, EN => n4987, Z 
                           => data_out_port_b(17));
   data_out_port_b_tri_18_inst : TBUF_X1 port map( A => n1791, EN => n4987, Z 
                           => data_out_port_b(18));
   data_out_port_b_tri_19_inst : TBUF_X1 port map( A => n1790, EN => n4987, Z 
                           => data_out_port_b(19));
   data_out_port_b_tri_20_inst : TBUF_X1 port map( A => n1789, EN => n4987, Z 
                           => data_out_port_b(20));
   data_out_port_b_tri_21_inst : TBUF_X1 port map( A => n1788, EN => n4987, Z 
                           => data_out_port_b(21));
   data_out_port_b_tri_22_inst : TBUF_X1 port map( A => n1787, EN => n4987, Z 
                           => data_out_port_b(22));
   data_out_port_b_tri_23_inst : TBUF_X1 port map( A => n1786, EN => n4987, Z 
                           => data_out_port_b(23));
   U3 : BUF_X1 port map( A => n555, Z => n4979);
   U4 : BUF_X1 port map( A => n555, Z => n4980);
   U5 : BUF_X1 port map( A => n1659, Z => n4886);
   U6 : BUF_X1 port map( A => n1659, Z => n4887);
   U7 : BUF_X1 port map( A => n555, Z => n4981);
   U8 : BUF_X1 port map( A => n1659, Z => n4888);
   U9 : BUF_X1 port map( A => n598, Z => n4907);
   U10 : BUF_X1 port map( A => n605, Z => n4895);
   U11 : BUF_X1 port map( A => n598, Z => n4908);
   U12 : BUF_X1 port map( A => n605, Z => n4896);
   U13 : BUF_X1 port map( A => n560, Z => n4973);
   U14 : BUF_X1 port map( A => n567, Z => n4961);
   U15 : BUF_X1 port map( A => n574, Z => n4949);
   U16 : BUF_X1 port map( A => n581, Z => n4937);
   U17 : BUF_X1 port map( A => n595, Z => n4916);
   U18 : BUF_X1 port map( A => n560, Z => n4974);
   U19 : BUF_X1 port map( A => n567, Z => n4962);
   U20 : BUF_X1 port map( A => n574, Z => n4950);
   U21 : BUF_X1 port map( A => n581, Z => n4938);
   U22 : BUF_X1 port map( A => n595, Z => n4917);
   U23 : BUF_X1 port map( A => n562, Z => n4967);
   U24 : BUF_X1 port map( A => n569, Z => n4955);
   U25 : BUF_X1 port map( A => n576, Z => n4943);
   U26 : BUF_X1 port map( A => n590, Z => n4922);
   U27 : BUF_X1 port map( A => n562, Z => n4968);
   U28 : BUF_X1 port map( A => n569, Z => n4956);
   U29 : BUF_X1 port map( A => n576, Z => n4944);
   U30 : BUF_X1 port map( A => n590, Z => n4923);
   U31 : BUF_X1 port map( A => n583, Z => n4931);
   U32 : BUF_X1 port map( A => n583, Z => n4932);
   U33 : BUF_X1 port map( A => n561, Z => n4970);
   U34 : BUF_X1 port map( A => n568, Z => n4958);
   U35 : BUF_X1 port map( A => n575, Z => n4946);
   U36 : BUF_X1 port map( A => n582, Z => n4934);
   U37 : BUF_X1 port map( A => n596, Z => n4913);
   U38 : BUF_X1 port map( A => n561, Z => n4971);
   U39 : BUF_X1 port map( A => n568, Z => n4959);
   U40 : BUF_X1 port map( A => n575, Z => n4947);
   U41 : BUF_X1 port map( A => n582, Z => n4935);
   U42 : BUF_X1 port map( A => n596, Z => n4914);
   U43 : BUF_X1 port map( A => n1692, Z => n4811);
   U44 : BUF_X1 port map( A => n1697, Z => n4799);
   U45 : BUF_X1 port map( A => n1682, Z => n4835);
   U46 : BUF_X1 port map( A => n1692, Z => n4812);
   U47 : BUF_X1 port map( A => n1697, Z => n4800);
   U48 : BUF_X1 port map( A => n1682, Z => n4836);
   U49 : BUF_X1 port map( A => n1693, Z => n4808);
   U50 : BUF_X1 port map( A => n1698, Z => n4796);
   U51 : BUF_X1 port map( A => n1683, Z => n4832);
   U52 : BUF_X1 port map( A => n1693, Z => n4809);
   U53 : BUF_X1 port map( A => n1698, Z => n4797);
   U54 : BUF_X1 port map( A => n1683, Z => n4833);
   U55 : BUF_X1 port map( A => n1660, Z => n4883);
   U56 : BUF_X1 port map( A => n1665, Z => n4871);
   U57 : BUF_X1 port map( A => n1670, Z => n4859);
   U58 : BUF_X1 port map( A => n1675, Z => n4847);
   U59 : BUF_X1 port map( A => n1685, Z => n4826);
   U60 : BUF_X1 port map( A => n1660, Z => n4884);
   U61 : BUF_X1 port map( A => n1665, Z => n4872);
   U62 : BUF_X1 port map( A => n1670, Z => n4860);
   U63 : BUF_X1 port map( A => n1675, Z => n4848);
   U64 : BUF_X1 port map( A => n1685, Z => n4827);
   U65 : BUF_X1 port map( A => n1689, Z => n4817);
   U66 : BUF_X1 port map( A => n1694, Z => n4805);
   U67 : BUF_X1 port map( A => n1689, Z => n4818);
   U68 : BUF_X1 port map( A => n1694, Z => n4806);
   U69 : BUF_X1 port map( A => n1679, Z => n4838);
   U70 : BUF_X1 port map( A => n1679, Z => n4839);
   U71 : BUF_X1 port map( A => n602, Z => n4901);
   U72 : BUF_X1 port map( A => n609, Z => n4889);
   U73 : BUF_X1 port map( A => n588, Z => n4925);
   U74 : BUF_X1 port map( A => n602, Z => n4902);
   U75 : BUF_X1 port map( A => n609, Z => n4890);
   U76 : BUF_X1 port map( A => n588, Z => n4926);
   U77 : BUF_X1 port map( A => n1662, Z => n4880);
   U78 : BUF_X1 port map( A => n1667, Z => n4868);
   U79 : BUF_X1 port map( A => n1672, Z => n4856);
   U80 : BUF_X1 port map( A => n1677, Z => n4844);
   U81 : BUF_X1 port map( A => n1687, Z => n4823);
   U82 : BUF_X1 port map( A => n1662, Z => n4881);
   U83 : BUF_X1 port map( A => n1667, Z => n4869);
   U84 : BUF_X1 port map( A => n1672, Z => n4857);
   U85 : BUF_X1 port map( A => n1677, Z => n4845);
   U86 : BUF_X1 port map( A => n1687, Z => n4824);
   U87 : BUF_X1 port map( A => n1690, Z => n4814);
   U88 : BUF_X1 port map( A => n1695, Z => n4802);
   U89 : BUF_X1 port map( A => n1690, Z => n4815);
   U90 : BUF_X1 port map( A => n1695, Z => n4803);
   U91 : BUF_X1 port map( A => n598, Z => n4909);
   U92 : BUF_X1 port map( A => n605, Z => n4897);
   U93 : BUF_X1 port map( A => n597, Z => n4910);
   U94 : BUF_X1 port map( A => n604, Z => n4898);
   U95 : BUF_X1 port map( A => n597, Z => n4911);
   U96 : BUF_X1 port map( A => n604, Z => n4899);
   U97 : BUF_X1 port map( A => n600, Z => n4904);
   U98 : BUF_X1 port map( A => n607, Z => n4892);
   U99 : BUF_X1 port map( A => n586, Z => n4928);
   U100 : BUF_X1 port map( A => n600, Z => n4905);
   U101 : BUF_X1 port map( A => n607, Z => n4893);
   U102 : BUF_X1 port map( A => n586, Z => n4929);
   U103 : BUF_X1 port map( A => n1664, Z => n4874);
   U104 : BUF_X1 port map( A => n1669, Z => n4862);
   U105 : BUF_X1 port map( A => n1674, Z => n4850);
   U106 : BUF_X1 port map( A => n1684, Z => n4829);
   U107 : BUF_X1 port map( A => n1664, Z => n4875);
   U108 : BUF_X1 port map( A => n1669, Z => n4863);
   U109 : BUF_X1 port map( A => n1674, Z => n4851);
   U110 : BUF_X1 port map( A => n1684, Z => n4830);
   U111 : BUF_X1 port map( A => n569, Z => n4957);
   U112 : BUF_X1 port map( A => n560, Z => n4975);
   U113 : BUF_X1 port map( A => n567, Z => n4963);
   U114 : BUF_X1 port map( A => n574, Z => n4951);
   U115 : BUF_X1 port map( A => n581, Z => n4939);
   U116 : BUF_X1 port map( A => n595, Z => n4918);
   U117 : BUF_X1 port map( A => n562, Z => n4969);
   U118 : BUF_X1 port map( A => n576, Z => n4945);
   U119 : BUF_X1 port map( A => n590, Z => n4924);
   U120 : BUF_X1 port map( A => n583, Z => n4933);
   U121 : BUF_X1 port map( A => n561, Z => n4972);
   U122 : BUF_X1 port map( A => n568, Z => n4960);
   U123 : BUF_X1 port map( A => n575, Z => n4948);
   U124 : BUF_X1 port map( A => n582, Z => n4936);
   U125 : BUF_X1 port map( A => n596, Z => n4915);
   U126 : BUF_X1 port map( A => n1692, Z => n4813);
   U127 : BUF_X1 port map( A => n1697, Z => n4801);
   U128 : BUF_X1 port map( A => n1682, Z => n4837);
   U129 : BUF_X1 port map( A => n557, Z => n4976);
   U130 : BUF_X1 port map( A => n564, Z => n4964);
   U131 : BUF_X1 port map( A => n571, Z => n4952);
   U132 : BUF_X1 port map( A => n578, Z => n4940);
   U133 : BUF_X1 port map( A => n592, Z => n4919);
   U134 : BUF_X1 port map( A => n557, Z => n4977);
   U135 : BUF_X1 port map( A => n564, Z => n4965);
   U136 : BUF_X1 port map( A => n571, Z => n4953);
   U137 : BUF_X1 port map( A => n578, Z => n4941);
   U138 : BUF_X1 port map( A => n592, Z => n4920);
   U139 : BUF_X1 port map( A => n1693, Z => n4810);
   U140 : BUF_X1 port map( A => n1698, Z => n4798);
   U141 : BUF_X1 port map( A => n1683, Z => n4834);
   U142 : BUF_X1 port map( A => n1663, Z => n4877);
   U143 : BUF_X1 port map( A => n1668, Z => n4865);
   U144 : BUF_X1 port map( A => n1673, Z => n4853);
   U145 : BUF_X1 port map( A => n1678, Z => n4841);
   U146 : BUF_X1 port map( A => n1688, Z => n4820);
   U147 : BUF_X1 port map( A => n1663, Z => n4878);
   U148 : BUF_X1 port map( A => n1668, Z => n4866);
   U149 : BUF_X1 port map( A => n1673, Z => n4854);
   U150 : BUF_X1 port map( A => n1678, Z => n4842);
   U151 : BUF_X1 port map( A => n1688, Z => n4821);
   U152 : BUF_X1 port map( A => n1660, Z => n4885);
   U153 : BUF_X1 port map( A => n1665, Z => n4873);
   U154 : BUF_X1 port map( A => n1670, Z => n4861);
   U155 : BUF_X1 port map( A => n1675, Z => n4849);
   U156 : BUF_X1 port map( A => n1685, Z => n4828);
   U157 : BUF_X1 port map( A => n1689, Z => n4819);
   U158 : BUF_X1 port map( A => n1694, Z => n4807);
   U159 : BUF_X1 port map( A => n1679, Z => n4840);
   U160 : BUF_X1 port map( A => n602, Z => n4903);
   U161 : BUF_X1 port map( A => n609, Z => n4891);
   U162 : BUF_X1 port map( A => n588, Z => n4927);
   U163 : BUF_X1 port map( A => n1662, Z => n4882);
   U164 : BUF_X1 port map( A => n1667, Z => n4870);
   U165 : BUF_X1 port map( A => n1672, Z => n4858);
   U166 : BUF_X1 port map( A => n1677, Z => n4846);
   U167 : BUF_X1 port map( A => n1687, Z => n4825);
   U168 : BUF_X1 port map( A => n1690, Z => n4816);
   U169 : BUF_X1 port map( A => n1695, Z => n4804);
   U170 : BUF_X1 port map( A => n597, Z => n4912);
   U171 : BUF_X1 port map( A => n604, Z => n4900);
   U172 : BUF_X1 port map( A => n600, Z => n4906);
   U173 : BUF_X1 port map( A => n607, Z => n4894);
   U174 : BUF_X1 port map( A => n586, Z => n4930);
   U175 : BUF_X1 port map( A => n1669, Z => n4864);
   U176 : BUF_X1 port map( A => n1674, Z => n4852);
   U177 : BUF_X1 port map( A => n1664, Z => n4876);
   U178 : BUF_X1 port map( A => n1684, Z => n4831);
   U179 : BUF_X1 port map( A => n592, Z => n4921);
   U180 : BUF_X1 port map( A => n557, Z => n4978);
   U181 : BUF_X1 port map( A => n564, Z => n4966);
   U182 : BUF_X1 port map( A => n571, Z => n4954);
   U183 : BUF_X1 port map( A => n578, Z => n4942);
   U184 : BUF_X1 port map( A => n1663, Z => n4879);
   U185 : BUF_X1 port map( A => n1668, Z => n4867);
   U186 : BUF_X1 port map( A => n1673, Z => n4855);
   U187 : BUF_X1 port map( A => n1678, Z => n4843);
   U188 : BUF_X1 port map( A => n1688, Z => n4822);
   U189 : NAND2_X1 port map( A1 => n2287, A2 => n2288, ZN => n1659);
   U190 : NAND2_X1 port map( A1 => n1617, A2 => n1618, ZN => n555);
   U191 : BUF_X1 port map( A => n2952, Z => n5105);
   U192 : BUF_X1 port map( A => n2952, Z => n5106);
   U193 : BUF_X1 port map( A => n2955, Z => n5102);
   U194 : BUF_X1 port map( A => n2955, Z => n5103);
   U195 : BUF_X1 port map( A => n2958, Z => n5099);
   U196 : BUF_X1 port map( A => n2958, Z => n5100);
   U197 : BUF_X1 port map( A => n2961, Z => n5096);
   U198 : BUF_X1 port map( A => n2961, Z => n5097);
   U199 : BUF_X1 port map( A => n2964, Z => n5093);
   U200 : BUF_X1 port map( A => n2964, Z => n5094);
   U201 : BUF_X1 port map( A => n2967, Z => n5090);
   U202 : BUF_X1 port map( A => n2967, Z => n5091);
   U203 : BUF_X1 port map( A => n2970, Z => n5087);
   U204 : BUF_X1 port map( A => n2970, Z => n5088);
   U205 : BUF_X1 port map( A => n2973, Z => n5084);
   U206 : BUF_X1 port map( A => n2973, Z => n5085);
   U207 : BUF_X1 port map( A => n2883, Z => n5174);
   U208 : BUF_X1 port map( A => n2883, Z => n5175);
   U209 : BUF_X1 port map( A => n2886, Z => n5171);
   U210 : BUF_X1 port map( A => n2886, Z => n5172);
   U211 : BUF_X1 port map( A => n2889, Z => n5168);
   U212 : BUF_X1 port map( A => n2889, Z => n5169);
   U213 : BUF_X1 port map( A => n2892, Z => n5165);
   U214 : BUF_X1 port map( A => n2892, Z => n5166);
   U215 : BUF_X1 port map( A => n2895, Z => n5162);
   U216 : BUF_X1 port map( A => n2895, Z => n5163);
   U217 : BUF_X1 port map( A => n2898, Z => n5159);
   U218 : BUF_X1 port map( A => n2898, Z => n5160);
   U219 : BUF_X1 port map( A => n2901, Z => n5156);
   U220 : BUF_X1 port map( A => n2901, Z => n5157);
   U221 : BUF_X1 port map( A => n2904, Z => n5153);
   U222 : BUF_X1 port map( A => n2904, Z => n5154);
   U223 : BUF_X1 port map( A => n2907, Z => n5150);
   U224 : BUF_X1 port map( A => n2907, Z => n5151);
   U225 : BUF_X1 port map( A => n2910, Z => n5147);
   U226 : BUF_X1 port map( A => n2910, Z => n5148);
   U227 : BUF_X1 port map( A => n2913, Z => n5144);
   U228 : BUF_X1 port map( A => n2913, Z => n5145);
   U229 : BUF_X1 port map( A => n2916, Z => n5141);
   U230 : BUF_X1 port map( A => n2916, Z => n5142);
   U231 : BUF_X1 port map( A => n2919, Z => n5138);
   U232 : BUF_X1 port map( A => n2919, Z => n5139);
   U233 : BUF_X1 port map( A => n2922, Z => n5135);
   U234 : BUF_X1 port map( A => n2922, Z => n5136);
   U235 : BUF_X1 port map( A => n2925, Z => n5132);
   U236 : BUF_X1 port map( A => n2925, Z => n5133);
   U237 : BUF_X1 port map( A => n2928, Z => n5129);
   U238 : BUF_X1 port map( A => n2928, Z => n5130);
   U239 : BUF_X1 port map( A => n2931, Z => n5126);
   U240 : BUF_X1 port map( A => n2931, Z => n5127);
   U241 : BUF_X1 port map( A => n2934, Z => n5123);
   U242 : BUF_X1 port map( A => n2934, Z => n5124);
   U243 : BUF_X1 port map( A => n2937, Z => n5120);
   U244 : BUF_X1 port map( A => n2937, Z => n5121);
   U245 : BUF_X1 port map( A => n2940, Z => n5117);
   U246 : BUF_X1 port map( A => n2940, Z => n5118);
   U247 : BUF_X1 port map( A => n2943, Z => n5114);
   U248 : BUF_X1 port map( A => n2943, Z => n5115);
   U249 : BUF_X1 port map( A => n2946, Z => n5111);
   U250 : BUF_X1 port map( A => n2946, Z => n5112);
   U251 : BUF_X1 port map( A => n2949, Z => n5108);
   U252 : BUF_X1 port map( A => n2949, Z => n5109);
   U253 : BUF_X1 port map( A => n2952, Z => n5107);
   U254 : BUF_X1 port map( A => n2955, Z => n5104);
   U255 : BUF_X1 port map( A => n2958, Z => n5101);
   U256 : BUF_X1 port map( A => n2961, Z => n5098);
   U257 : BUF_X1 port map( A => n2964, Z => n5095);
   U258 : BUF_X1 port map( A => n2967, Z => n5092);
   U259 : BUF_X1 port map( A => n2970, Z => n5089);
   U260 : BUF_X1 port map( A => n2973, Z => n5086);
   U261 : BUF_X1 port map( A => n2883, Z => n5176);
   U262 : BUF_X1 port map( A => n2886, Z => n5173);
   U263 : BUF_X1 port map( A => n2889, Z => n5170);
   U264 : BUF_X1 port map( A => n2892, Z => n5167);
   U265 : BUF_X1 port map( A => n2895, Z => n5164);
   U266 : BUF_X1 port map( A => n2898, Z => n5161);
   U267 : BUF_X1 port map( A => n2901, Z => n5158);
   U268 : BUF_X1 port map( A => n2904, Z => n5155);
   U269 : BUF_X1 port map( A => n2907, Z => n5152);
   U270 : BUF_X1 port map( A => n2910, Z => n5149);
   U271 : BUF_X1 port map( A => n2913, Z => n5146);
   U272 : BUF_X1 port map( A => n2916, Z => n5143);
   U273 : BUF_X1 port map( A => n2919, Z => n5140);
   U274 : BUF_X1 port map( A => n2922, Z => n5137);
   U275 : BUF_X1 port map( A => n2925, Z => n5134);
   U276 : BUF_X1 port map( A => n2928, Z => n5131);
   U277 : BUF_X1 port map( A => n2931, Z => n5128);
   U278 : BUF_X1 port map( A => n2934, Z => n5125);
   U279 : BUF_X1 port map( A => n2937, Z => n5122);
   U280 : BUF_X1 port map( A => n2940, Z => n5119);
   U281 : BUF_X1 port map( A => n2943, Z => n5116);
   U282 : BUF_X1 port map( A => n2946, Z => n5113);
   U283 : BUF_X1 port map( A => n2949, Z => n5110);
   U284 : NOR2_X1 port map( A1 => n2305, A2 => n2306, ZN => n2287);
   U285 : NOR2_X1 port map( A1 => n1649, A2 => n1650, ZN => n1617);
   U286 : NOR3_X1 port map( A1 => n1637, A2 => n1641, A3 => n1642, ZN => n1618)
                           ;
   U287 : NOR3_X1 port map( A1 => n2299, A2 => n2301, A3 => n2302, ZN => n2288)
                           ;
   U288 : NOR4_X1 port map( A1 => n2005, A2 => n2006, A3 => n2007, A4 => n2008,
                           ZN => n2004);
   U289 : OAI221_X1 port map( B1 => n1090, B2 => n4851, C1 => n1091, C2 => 
                           n4848, A => n2012, ZN => n2005);
   U290 : OAI221_X1 port map( B1 => n1087, B2 => n4863, C1 => n1088, C2 => 
                           n4860, A => n2011, ZN => n2006);
   U291 : OAI221_X1 port map( B1 => n1084, B2 => n4875, C1 => n1085, C2 => 
                           n4872, A => n2010, ZN => n2007);
   U292 : NOR4_X1 port map( A1 => n1988, A2 => n1989, A3 => n1990, A4 => n1991,
                           ZN => n1987);
   U293 : OAI221_X1 port map( B1 => n1057, B2 => n4851, C1 => n1058, C2 => 
                           n4848, A => n1995, ZN => n1988);
   U294 : OAI221_X1 port map( B1 => n1054, B2 => n4863, C1 => n1055, C2 => 
                           n4860, A => n1994, ZN => n1989);
   U295 : OAI221_X1 port map( B1 => n1051, B2 => n4875, C1 => n1052, C2 => 
                           n4872, A => n1993, ZN => n1990);
   U296 : NOR4_X1 port map( A1 => n1971, A2 => n1972, A3 => n1973, A4 => n1974,
                           ZN => n1970);
   U297 : OAI221_X1 port map( B1 => n1024, B2 => n4851, C1 => n1025, C2 => 
                           n4848, A => n1978, ZN => n1971);
   U298 : OAI221_X1 port map( B1 => n1021, B2 => n4863, C1 => n1022, C2 => 
                           n4860, A => n1977, ZN => n1972);
   U299 : OAI221_X1 port map( B1 => n1018, B2 => n4875, C1 => n1019, C2 => 
                           n4872, A => n1976, ZN => n1973);
   U300 : NOR4_X1 port map( A1 => n1954, A2 => n1955, A3 => n1956, A4 => n1957,
                           ZN => n1953);
   U301 : OAI221_X1 port map( B1 => n991, B2 => n4851, C1 => n992, C2 => n4848,
                           A => n1961, ZN => n1954);
   U302 : OAI221_X1 port map( B1 => n988, B2 => n4863, C1 => n989, C2 => n4860,
                           A => n1960, ZN => n1955);
   U303 : OAI221_X1 port map( B1 => n985, B2 => n4875, C1 => n986, C2 => n4872,
                           A => n1959, ZN => n1956);
   U304 : NOR4_X1 port map( A1 => n1937, A2 => n1938, A3 => n1939, A4 => n1940,
                           ZN => n1936);
   U305 : OAI221_X1 port map( B1 => n958, B2 => n4851, C1 => n959, C2 => n4848,
                           A => n1944, ZN => n1937);
   U306 : OAI221_X1 port map( B1 => n955, B2 => n4863, C1 => n956, C2 => n4860,
                           A => n1943, ZN => n1938);
   U307 : OAI221_X1 port map( B1 => n952, B2 => n4875, C1 => n953, C2 => n4872,
                           A => n1942, ZN => n1939);
   U308 : NOR4_X1 port map( A1 => n1920, A2 => n1921, A3 => n1922, A4 => n1923,
                           ZN => n1919);
   U309 : OAI221_X1 port map( B1 => n925, B2 => n4851, C1 => n926, C2 => n4848,
                           A => n1927, ZN => n1920);
   U310 : OAI221_X1 port map( B1 => n922, B2 => n4863, C1 => n923, C2 => n4860,
                           A => n1926, ZN => n1921);
   U311 : OAI221_X1 port map( B1 => n919, B2 => n4875, C1 => n920, C2 => n4872,
                           A => n1925, ZN => n1922);
   U312 : NOR4_X1 port map( A1 => n1903, A2 => n1904, A3 => n1905, A4 => n1906,
                           ZN => n1902);
   U313 : OAI221_X1 port map( B1 => n892, B2 => n4851, C1 => n893, C2 => n4848,
                           A => n1910, ZN => n1903);
   U314 : OAI221_X1 port map( B1 => n889, B2 => n4863, C1 => n890, C2 => n4860,
                           A => n1909, ZN => n1904);
   U315 : OAI221_X1 port map( B1 => n886, B2 => n4875, C1 => n887, C2 => n4872,
                           A => n1908, ZN => n1905);
   U316 : NOR4_X1 port map( A1 => n1886, A2 => n1887, A3 => n1888, A4 => n1889,
                           ZN => n1885);
   U317 : OAI221_X1 port map( B1 => n859, B2 => n4851, C1 => n860, C2 => n4848,
                           A => n1893, ZN => n1886);
   U318 : OAI221_X1 port map( B1 => n856, B2 => n4863, C1 => n857, C2 => n4860,
                           A => n1892, ZN => n1887);
   U319 : OAI221_X1 port map( B1 => n853, B2 => n4875, C1 => n854, C2 => n4872,
                           A => n1891, ZN => n1888);
   U320 : NOR4_X1 port map( A1 => n2277, A2 => n2278, A3 => n2279, A4 => n2280,
                           ZN => n2276);
   U321 : OAI221_X1 port map( B1 => n1630, B2 => n4850, C1 => n1631, C2 => 
                           n4847, A => n2296, ZN => n2277);
   U322 : OAI221_X1 port map( B1 => n1625, B2 => n4862, C1 => n1626, C2 => 
                           n4859, A => n2293, ZN => n2278);
   U323 : OAI221_X1 port map( B1 => n1619, B2 => n4874, C1 => n1620, C2 => 
                           n4871, A => n2289, ZN => n2279);
   U324 : NOR4_X1 port map( A1 => n2260, A2 => n2261, A3 => n2262, A4 => n2263,
                           ZN => n2259);
   U325 : OAI221_X1 port map( B1 => n1585, B2 => n4850, C1 => n1586, C2 => 
                           n4847, A => n2267, ZN => n2260);
   U326 : OAI221_X1 port map( B1 => n1582, B2 => n4862, C1 => n1583, C2 => 
                           n4859, A => n2266, ZN => n2261);
   U327 : OAI221_X1 port map( B1 => n1579, B2 => n4874, C1 => n1580, C2 => 
                           n4871, A => n2265, ZN => n2262);
   U328 : NOR4_X1 port map( A1 => n2243, A2 => n2244, A3 => n2245, A4 => n2246,
                           ZN => n2242);
   U329 : OAI221_X1 port map( B1 => n1552, B2 => n4850, C1 => n1553, C2 => 
                           n4847, A => n2250, ZN => n2243);
   U330 : OAI221_X1 port map( B1 => n1549, B2 => n4862, C1 => n1550, C2 => 
                           n4859, A => n2249, ZN => n2244);
   U331 : OAI221_X1 port map( B1 => n1546, B2 => n4874, C1 => n1547, C2 => 
                           n4871, A => n2248, ZN => n2245);
   U332 : NOR4_X1 port map( A1 => n2226, A2 => n2227, A3 => n2228, A4 => n2229,
                           ZN => n2225);
   U333 : OAI221_X1 port map( B1 => n1519, B2 => n4850, C1 => n1520, C2 => 
                           n4847, A => n2233, ZN => n2226);
   U334 : OAI221_X1 port map( B1 => n1516, B2 => n4862, C1 => n1517, C2 => 
                           n4859, A => n2232, ZN => n2227);
   U335 : OAI221_X1 port map( B1 => n1513, B2 => n4874, C1 => n1514, C2 => 
                           n4871, A => n2231, ZN => n2228);
   U336 : NOR4_X1 port map( A1 => n2209, A2 => n2210, A3 => n2211, A4 => n2212,
                           ZN => n2208);
   U337 : OAI221_X1 port map( B1 => n1486, B2 => n4850, C1 => n1487, C2 => 
                           n4847, A => n2216, ZN => n2209);
   U338 : OAI221_X1 port map( B1 => n1483, B2 => n4862, C1 => n1484, C2 => 
                           n4859, A => n2215, ZN => n2210);
   U339 : OAI221_X1 port map( B1 => n1480, B2 => n4874, C1 => n1481, C2 => 
                           n4871, A => n2214, ZN => n2211);
   U340 : NOR4_X1 port map( A1 => n2192, A2 => n2193, A3 => n2194, A4 => n2195,
                           ZN => n2191);
   U341 : OAI221_X1 port map( B1 => n1453, B2 => n4850, C1 => n1454, C2 => 
                           n4847, A => n2199, ZN => n2192);
   U342 : OAI221_X1 port map( B1 => n1450, B2 => n4862, C1 => n1451, C2 => 
                           n4859, A => n2198, ZN => n2193);
   U343 : OAI221_X1 port map( B1 => n1447, B2 => n4874, C1 => n1448, C2 => 
                           n4871, A => n2197, ZN => n2194);
   U344 : NOR4_X1 port map( A1 => n2175, A2 => n2176, A3 => n2177, A4 => n2178,
                           ZN => n2174);
   U345 : OAI221_X1 port map( B1 => n1420, B2 => n4850, C1 => n1421, C2 => 
                           n4847, A => n2182, ZN => n2175);
   U346 : OAI221_X1 port map( B1 => n1417, B2 => n4862, C1 => n1418, C2 => 
                           n4859, A => n2181, ZN => n2176);
   U347 : OAI221_X1 port map( B1 => n1414, B2 => n4874, C1 => n1415, C2 => 
                           n4871, A => n2180, ZN => n2177);
   U348 : NOR4_X1 port map( A1 => n2158, A2 => n2159, A3 => n2160, A4 => n2161,
                           ZN => n2157);
   U349 : OAI221_X1 port map( B1 => n1387, B2 => n4850, C1 => n1388, C2 => 
                           n4847, A => n2165, ZN => n2158);
   U350 : OAI221_X1 port map( B1 => n1384, B2 => n4862, C1 => n1385, C2 => 
                           n4859, A => n2164, ZN => n2159);
   U351 : OAI221_X1 port map( B1 => n1381, B2 => n4874, C1 => n1382, C2 => 
                           n4871, A => n2163, ZN => n2160);
   U352 : NOR4_X1 port map( A1 => n2141, A2 => n2142, A3 => n2143, A4 => n2144,
                           ZN => n2140);
   U353 : OAI221_X1 port map( B1 => n1354, B2 => n4850, C1 => n1355, C2 => 
                           n4847, A => n2148, ZN => n2141);
   U354 : OAI221_X1 port map( B1 => n1351, B2 => n4862, C1 => n1352, C2 => 
                           n4859, A => n2147, ZN => n2142);
   U355 : OAI221_X1 port map( B1 => n1348, B2 => n4874, C1 => n1349, C2 => 
                           n4871, A => n2146, ZN => n2143);
   U356 : NOR4_X1 port map( A1 => n2124, A2 => n2125, A3 => n2126, A4 => n2127,
                           ZN => n2123);
   U357 : OAI221_X1 port map( B1 => n1321, B2 => n4850, C1 => n1322, C2 => 
                           n4847, A => n2131, ZN => n2124);
   U358 : OAI221_X1 port map( B1 => n1318, B2 => n4862, C1 => n1319, C2 => 
                           n4859, A => n2130, ZN => n2125);
   U359 : OAI221_X1 port map( B1 => n1315, B2 => n4874, C1 => n1316, C2 => 
                           n4871, A => n2129, ZN => n2126);
   U360 : NOR4_X1 port map( A1 => n2107, A2 => n2108, A3 => n2109, A4 => n2110,
                           ZN => n2106);
   U361 : OAI221_X1 port map( B1 => n1288, B2 => n4850, C1 => n1289, C2 => 
                           n4847, A => n2114, ZN => n2107);
   U362 : OAI221_X1 port map( B1 => n1285, B2 => n4862, C1 => n1286, C2 => 
                           n4859, A => n2113, ZN => n2108);
   U363 : OAI221_X1 port map( B1 => n1282, B2 => n4874, C1 => n1283, C2 => 
                           n4871, A => n2112, ZN => n2109);
   U364 : NOR4_X1 port map( A1 => n2090, A2 => n2091, A3 => n2092, A4 => n2093,
                           ZN => n2089);
   U365 : OAI221_X1 port map( B1 => n1255, B2 => n4850, C1 => n1256, C2 => 
                           n4847, A => n2097, ZN => n2090);
   U366 : OAI221_X1 port map( B1 => n1252, B2 => n4862, C1 => n1253, C2 => 
                           n4859, A => n2096, ZN => n2091);
   U367 : OAI221_X1 port map( B1 => n1249, B2 => n4874, C1 => n1250, C2 => 
                           n4871, A => n2095, ZN => n2092);
   U368 : NOR4_X1 port map( A1 => n2073, A2 => n2074, A3 => n2075, A4 => n2076,
                           ZN => n2072);
   U369 : OAI221_X1 port map( B1 => n1222, B2 => n4851, C1 => n1223, C2 => 
                           n4848, A => n2080, ZN => n2073);
   U370 : OAI221_X1 port map( B1 => n1219, B2 => n4863, C1 => n1220, C2 => 
                           n4860, A => n2079, ZN => n2074);
   U371 : OAI221_X1 port map( B1 => n1216, B2 => n4875, C1 => n1217, C2 => 
                           n4872, A => n2078, ZN => n2075);
   U372 : NOR4_X1 port map( A1 => n2056, A2 => n2057, A3 => n2058, A4 => n2059,
                           ZN => n2055);
   U373 : OAI221_X1 port map( B1 => n1189, B2 => n4851, C1 => n1190, C2 => 
                           n4848, A => n2063, ZN => n2056);
   U374 : OAI221_X1 port map( B1 => n1186, B2 => n4863, C1 => n1187, C2 => 
                           n4860, A => n2062, ZN => n2057);
   U375 : OAI221_X1 port map( B1 => n1183, B2 => n4875, C1 => n1184, C2 => 
                           n4872, A => n2061, ZN => n2058);
   U376 : NOR4_X1 port map( A1 => n2039, A2 => n2040, A3 => n2041, A4 => n2042,
                           ZN => n2038);
   U377 : OAI221_X1 port map( B1 => n1156, B2 => n4851, C1 => n1157, C2 => 
                           n4848, A => n2046, ZN => n2039);
   U378 : OAI221_X1 port map( B1 => n1153, B2 => n4863, C1 => n1154, C2 => 
                           n4860, A => n2045, ZN => n2040);
   U379 : OAI221_X1 port map( B1 => n1150, B2 => n4875, C1 => n1151, C2 => 
                           n4872, A => n2044, ZN => n2041);
   U380 : NOR4_X1 port map( A1 => n2022, A2 => n2023, A3 => n2024, A4 => n2025,
                           ZN => n2021);
   U381 : OAI221_X1 port map( B1 => n1123, B2 => n4851, C1 => n1124, C2 => 
                           n4848, A => n2029, ZN => n2022);
   U382 : OAI221_X1 port map( B1 => n1120, B2 => n4863, C1 => n1121, C2 => 
                           n4860, A => n2028, ZN => n2023);
   U383 : OAI221_X1 port map( B1 => n1117, B2 => n4875, C1 => n1118, C2 => 
                           n4872, A => n2027, ZN => n2024);
   U384 : NOR4_X1 port map( A1 => n1869, A2 => n1870, A3 => n1871, A4 => n1872,
                           ZN => n1868);
   U385 : OAI221_X1 port map( B1 => n826, B2 => n4852, C1 => n827, C2 => n4849,
                           A => n1876, ZN => n1869);
   U386 : OAI221_X1 port map( B1 => n823, B2 => n4864, C1 => n824, C2 => n4861,
                           A => n1875, ZN => n1870);
   U387 : OAI221_X1 port map( B1 => n820, B2 => n4876, C1 => n821, C2 => n4873,
                           A => n1874, ZN => n1871);
   U388 : NOR4_X1 port map( A1 => n1852, A2 => n1853, A3 => n1854, A4 => n1855,
                           ZN => n1851);
   U389 : OAI221_X1 port map( B1 => n793, B2 => n4852, C1 => n794, C2 => n4849,
                           A => n1859, ZN => n1852);
   U390 : OAI221_X1 port map( B1 => n790, B2 => n4864, C1 => n791, C2 => n4861,
                           A => n1858, ZN => n1853);
   U391 : OAI221_X1 port map( B1 => n787, B2 => n4876, C1 => n788, C2 => n4873,
                           A => n1857, ZN => n1854);
   U392 : NOR4_X1 port map( A1 => n1771, A2 => n1772, A3 => n1773, A4 => n1774,
                           ZN => n1770);
   U393 : OAI221_X1 port map( B1 => n760, B2 => n4852, C1 => n761, C2 => n4849,
                           A => n1801, ZN => n1771);
   U394 : OAI221_X1 port map( B1 => n757, B2 => n4864, C1 => n758, C2 => n4861,
                           A => n1777, ZN => n1772);
   U395 : OAI221_X1 port map( B1 => n754, B2 => n4876, C1 => n755, C2 => n4873,
                           A => n1776, ZN => n1773);
   U396 : NOR4_X1 port map( A1 => n1754, A2 => n1755, A3 => n1756, A4 => n1757,
                           ZN => n1753);
   U397 : OAI221_X1 port map( B1 => n727, B2 => n4852, C1 => n728, C2 => n4849,
                           A => n1761, ZN => n1754);
   U398 : OAI221_X1 port map( B1 => n724, B2 => n4864, C1 => n725, C2 => n4861,
                           A => n1760, ZN => n1755);
   U399 : OAI221_X1 port map( B1 => n721, B2 => n4876, C1 => n722, C2 => n4873,
                           A => n1759, ZN => n1756);
   U400 : NOR4_X1 port map( A1 => n1737, A2 => n1738, A3 => n1739, A4 => n1740,
                           ZN => n1736);
   U401 : OAI221_X1 port map( B1 => n694, B2 => n4852, C1 => n695, C2 => n4849,
                           A => n1744, ZN => n1737);
   U402 : OAI221_X1 port map( B1 => n691, B2 => n4864, C1 => n692, C2 => n4861,
                           A => n1743, ZN => n1738);
   U403 : OAI221_X1 port map( B1 => n688, B2 => n4876, C1 => n689, C2 => n4873,
                           A => n1742, ZN => n1739);
   U404 : NOR4_X1 port map( A1 => n1720, A2 => n1721, A3 => n1722, A4 => n1723,
                           ZN => n1719);
   U405 : OAI221_X1 port map( B1 => n661, B2 => n4852, C1 => n662, C2 => n4849,
                           A => n1727, ZN => n1720);
   U406 : OAI221_X1 port map( B1 => n658, B2 => n4864, C1 => n659, C2 => n4861,
                           A => n1726, ZN => n1721);
   U407 : OAI221_X1 port map( B1 => n655, B2 => n4876, C1 => n656, C2 => n4873,
                           A => n1725, ZN => n1722);
   U408 : NOR4_X1 port map( A1 => n1703, A2 => n1704, A3 => n1705, A4 => n1706,
                           ZN => n1702);
   U409 : OAI221_X1 port map( B1 => n628, B2 => n4852, C1 => n629, C2 => n4849,
                           A => n1710, ZN => n1703);
   U410 : OAI221_X1 port map( B1 => n625, B2 => n4864, C1 => n626, C2 => n4861,
                           A => n1709, ZN => n1704);
   U411 : OAI221_X1 port map( B1 => n622, B2 => n4876, C1 => n623, C2 => n4873,
                           A => n1708, ZN => n1705);
   U412 : NOR4_X1 port map( A1 => n1655, A2 => n1656, A3 => n1657, A4 => n1658,
                           ZN => n1654);
   U413 : OAI221_X1 port map( B1 => n577, B2 => n4852, C1 => n579, C2 => n4849,
                           A => n1676, ZN => n1655);
   U414 : OAI221_X1 port map( B1 => n570, B2 => n4864, C1 => n572, C2 => n4861,
                           A => n1671, ZN => n1656);
   U415 : OAI221_X1 port map( B1 => n563, B2 => n4876, C1 => n565, C2 => n4873,
                           A => n1666, ZN => n1657);
   U416 : NOR4_X1 port map( A1 => n1077, A2 => n1078, A3 => n1079, A4 => n1080,
                           ZN => n1076);
   U417 : OAI221_X1 port map( B1 => n4944, B2 => n1090, C1 => n4941, C2 => 
                           n1091, A => n1092, ZN => n1077);
   U418 : OAI221_X1 port map( B1 => n4956, B2 => n1087, C1 => n4953, C2 => 
                           n1088, A => n1089, ZN => n1078);
   U419 : OAI221_X1 port map( B1 => n4968, B2 => n1084, C1 => n4965, C2 => 
                           n1085, A => n1086, ZN => n1079);
   U420 : NOR4_X1 port map( A1 => n1044, A2 => n1045, A3 => n1046, A4 => n1047,
                           ZN => n1043);
   U421 : OAI221_X1 port map( B1 => n4944, B2 => n1057, C1 => n4941, C2 => 
                           n1058, A => n1059, ZN => n1044);
   U422 : OAI221_X1 port map( B1 => n4956, B2 => n1054, C1 => n4953, C2 => 
                           n1055, A => n1056, ZN => n1045);
   U423 : OAI221_X1 port map( B1 => n4968, B2 => n1051, C1 => n4965, C2 => 
                           n1052, A => n1053, ZN => n1046);
   U424 : NOR4_X1 port map( A1 => n1011, A2 => n1012, A3 => n1013, A4 => n1014,
                           ZN => n1010);
   U425 : OAI221_X1 port map( B1 => n4944, B2 => n1024, C1 => n4941, C2 => 
                           n1025, A => n1026, ZN => n1011);
   U426 : OAI221_X1 port map( B1 => n4956, B2 => n1021, C1 => n4953, C2 => 
                           n1022, A => n1023, ZN => n1012);
   U427 : OAI221_X1 port map( B1 => n4968, B2 => n1018, C1 => n4965, C2 => 
                           n1019, A => n1020, ZN => n1013);
   U428 : NOR4_X1 port map( A1 => n978, A2 => n979, A3 => n980, A4 => n981, ZN 
                           => n977);
   U429 : OAI221_X1 port map( B1 => n4944, B2 => n991, C1 => n4941, C2 => n992,
                           A => n993, ZN => n978);
   U430 : OAI221_X1 port map( B1 => n4956, B2 => n988, C1 => n4953, C2 => n989,
                           A => n990, ZN => n979);
   U431 : OAI221_X1 port map( B1 => n4968, B2 => n985, C1 => n4965, C2 => n986,
                           A => n987, ZN => n980);
   U432 : NOR4_X1 port map( A1 => n945, A2 => n946, A3 => n947, A4 => n948, ZN 
                           => n944);
   U433 : OAI221_X1 port map( B1 => n4944, B2 => n958, C1 => n4941, C2 => n959,
                           A => n960, ZN => n945);
   U434 : OAI221_X1 port map( B1 => n4956, B2 => n955, C1 => n4953, C2 => n956,
                           A => n957, ZN => n946);
   U435 : OAI221_X1 port map( B1 => n4968, B2 => n952, C1 => n4965, C2 => n953,
                           A => n954, ZN => n947);
   U436 : NOR4_X1 port map( A1 => n912, A2 => n913, A3 => n914, A4 => n915, ZN 
                           => n911);
   U437 : OAI221_X1 port map( B1 => n4944, B2 => n925, C1 => n4941, C2 => n926,
                           A => n927, ZN => n912);
   U438 : OAI221_X1 port map( B1 => n4956, B2 => n922, C1 => n4953, C2 => n923,
                           A => n924, ZN => n913);
   U439 : OAI221_X1 port map( B1 => n4968, B2 => n919, C1 => n4965, C2 => n920,
                           A => n921, ZN => n914);
   U440 : NOR4_X1 port map( A1 => n879, A2 => n880, A3 => n881, A4 => n882, ZN 
                           => n878);
   U441 : OAI221_X1 port map( B1 => n4944, B2 => n892, C1 => n4941, C2 => n893,
                           A => n894, ZN => n879);
   U442 : OAI221_X1 port map( B1 => n4956, B2 => n889, C1 => n4953, C2 => n890,
                           A => n891, ZN => n880);
   U443 : OAI221_X1 port map( B1 => n4968, B2 => n886, C1 => n4965, C2 => n887,
                           A => n888, ZN => n881);
   U444 : NOR4_X1 port map( A1 => n846, A2 => n847, A3 => n848, A4 => n849, ZN 
                           => n845);
   U445 : OAI221_X1 port map( B1 => n4944, B2 => n859, C1 => n4941, C2 => n860,
                           A => n861, ZN => n846);
   U446 : OAI221_X1 port map( B1 => n4956, B2 => n856, C1 => n4953, C2 => n857,
                           A => n858, ZN => n847);
   U447 : OAI221_X1 port map( B1 => n4968, B2 => n853, C1 => n4965, C2 => n854,
                           A => n855, ZN => n848);
   U448 : NOR4_X1 port map( A1 => n813, A2 => n814, A3 => n815, A4 => n816, ZN 
                           => n812);
   U449 : OAI221_X1 port map( B1 => n4945, B2 => n826, C1 => n4942, C2 => n827,
                           A => n828, ZN => n813);
   U450 : OAI221_X1 port map( B1 => n4957, B2 => n823, C1 => n4954, C2 => n824,
                           A => n825, ZN => n814);
   U451 : OAI221_X1 port map( B1 => n4969, B2 => n820, C1 => n4966, C2 => n821,
                           A => n822, ZN => n815);
   U452 : NOR4_X1 port map( A1 => n780, A2 => n781, A3 => n782, A4 => n783, ZN 
                           => n779);
   U453 : OAI221_X1 port map( B1 => n4945, B2 => n793, C1 => n4942, C2 => n794,
                           A => n795, ZN => n780);
   U454 : OAI221_X1 port map( B1 => n4957, B2 => n790, C1 => n4954, C2 => n791,
                           A => n792, ZN => n781);
   U455 : OAI221_X1 port map( B1 => n4969, B2 => n787, C1 => n4966, C2 => n788,
                           A => n789, ZN => n782);
   U456 : NOR4_X1 port map( A1 => n747, A2 => n748, A3 => n749, A4 => n750, ZN 
                           => n746);
   U457 : OAI221_X1 port map( B1 => n4945, B2 => n760, C1 => n4942, C2 => n761,
                           A => n762, ZN => n747);
   U458 : OAI221_X1 port map( B1 => n4957, B2 => n757, C1 => n4954, C2 => n758,
                           A => n759, ZN => n748);
   U459 : OAI221_X1 port map( B1 => n4969, B2 => n754, C1 => n4966, C2 => n755,
                           A => n756, ZN => n749);
   U460 : NOR4_X1 port map( A1 => n714, A2 => n715, A3 => n716, A4 => n717, ZN 
                           => n713);
   U461 : OAI221_X1 port map( B1 => n4945, B2 => n727, C1 => n4942, C2 => n728,
                           A => n729, ZN => n714);
   U462 : OAI221_X1 port map( B1 => n4957, B2 => n724, C1 => n4954, C2 => n725,
                           A => n726, ZN => n715);
   U463 : OAI221_X1 port map( B1 => n4969, B2 => n721, C1 => n4966, C2 => n722,
                           A => n723, ZN => n716);
   U464 : NOR4_X1 port map( A1 => n681, A2 => n682, A3 => n683, A4 => n684, ZN 
                           => n680);
   U465 : OAI221_X1 port map( B1 => n4945, B2 => n694, C1 => n4942, C2 => n695,
                           A => n696, ZN => n681);
   U466 : OAI221_X1 port map( B1 => n4957, B2 => n691, C1 => n4954, C2 => n692,
                           A => n693, ZN => n682);
   U467 : OAI221_X1 port map( B1 => n4969, B2 => n688, C1 => n4966, C2 => n689,
                           A => n690, ZN => n683);
   U468 : NOR4_X1 port map( A1 => n648, A2 => n649, A3 => n650, A4 => n651, ZN 
                           => n647);
   U469 : OAI221_X1 port map( B1 => n4945, B2 => n661, C1 => n4942, C2 => n662,
                           A => n663, ZN => n648);
   U470 : OAI221_X1 port map( B1 => n4957, B2 => n658, C1 => n4954, C2 => n659,
                           A => n660, ZN => n649);
   U471 : OAI221_X1 port map( B1 => n4969, B2 => n655, C1 => n4966, C2 => n656,
                           A => n657, ZN => n650);
   U472 : NOR4_X1 port map( A1 => n615, A2 => n616, A3 => n617, A4 => n618, ZN 
                           => n614);
   U473 : OAI221_X1 port map( B1 => n4945, B2 => n628, C1 => n4942, C2 => n629,
                           A => n630, ZN => n615);
   U474 : OAI221_X1 port map( B1 => n4957, B2 => n625, C1 => n4954, C2 => n626,
                           A => n627, ZN => n616);
   U475 : OAI221_X1 port map( B1 => n4969, B2 => n622, C1 => n4966, C2 => n623,
                           A => n624, ZN => n617);
   U476 : NOR4_X1 port map( A1 => n551, A2 => n552, A3 => n553, A4 => n554, ZN 
                           => n550);
   U477 : OAI221_X1 port map( B1 => n4945, B2 => n577, C1 => n4942, C2 => n579,
                           A => n580, ZN => n551);
   U478 : OAI221_X1 port map( B1 => n4957, B2 => n570, C1 => n4954, C2 => n572,
                           A => n573, ZN => n552);
   U479 : OAI221_X1 port map( B1 => n4969, B2 => n563, C1 => n4966, C2 => n565,
                           A => n566, ZN => n553);
   U480 : NOR4_X1 port map( A1 => n1605, A2 => n1606, A3 => n1607, A4 => n1608,
                           ZN => n1604);
   U481 : OAI221_X1 port map( B1 => n4943, B2 => n1630, C1 => n4940, C2 => 
                           n1631, A => n1632, ZN => n1605);
   U482 : OAI221_X1 port map( B1 => n4955, B2 => n1625, C1 => n4952, C2 => 
                           n1626, A => n1627, ZN => n1606);
   U483 : OAI221_X1 port map( B1 => n4967, B2 => n1619, C1 => n4964, C2 => 
                           n1620, A => n1621, ZN => n1607);
   U484 : NOR4_X1 port map( A1 => n1572, A2 => n1573, A3 => n1574, A4 => n1575,
                           ZN => n1571);
   U485 : OAI221_X1 port map( B1 => n4943, B2 => n1585, C1 => n4940, C2 => 
                           n1586, A => n1587, ZN => n1572);
   U486 : OAI221_X1 port map( B1 => n4955, B2 => n1582, C1 => n4952, C2 => 
                           n1583, A => n1584, ZN => n1573);
   U487 : OAI221_X1 port map( B1 => n4967, B2 => n1579, C1 => n4964, C2 => 
                           n1580, A => n1581, ZN => n1574);
   U488 : NOR4_X1 port map( A1 => n1539, A2 => n1540, A3 => n1541, A4 => n1542,
                           ZN => n1538);
   U489 : OAI221_X1 port map( B1 => n4943, B2 => n1552, C1 => n4940, C2 => 
                           n1553, A => n1554, ZN => n1539);
   U490 : OAI221_X1 port map( B1 => n4955, B2 => n1549, C1 => n4952, C2 => 
                           n1550, A => n1551, ZN => n1540);
   U491 : OAI221_X1 port map( B1 => n4967, B2 => n1546, C1 => n4964, C2 => 
                           n1547, A => n1548, ZN => n1541);
   U492 : NOR4_X1 port map( A1 => n1506, A2 => n1507, A3 => n1508, A4 => n1509,
                           ZN => n1505);
   U493 : OAI221_X1 port map( B1 => n4943, B2 => n1519, C1 => n4940, C2 => 
                           n1520, A => n1521, ZN => n1506);
   U494 : OAI221_X1 port map( B1 => n4955, B2 => n1516, C1 => n4952, C2 => 
                           n1517, A => n1518, ZN => n1507);
   U495 : OAI221_X1 port map( B1 => n4967, B2 => n1513, C1 => n4964, C2 => 
                           n1514, A => n1515, ZN => n1508);
   U496 : NOR4_X1 port map( A1 => n1473, A2 => n1474, A3 => n1475, A4 => n1476,
                           ZN => n1472);
   U497 : OAI221_X1 port map( B1 => n4943, B2 => n1486, C1 => n4940, C2 => 
                           n1487, A => n1488, ZN => n1473);
   U498 : OAI221_X1 port map( B1 => n4955, B2 => n1483, C1 => n4952, C2 => 
                           n1484, A => n1485, ZN => n1474);
   U499 : OAI221_X1 port map( B1 => n4967, B2 => n1480, C1 => n4964, C2 => 
                           n1481, A => n1482, ZN => n1475);
   U500 : NOR4_X1 port map( A1 => n1440, A2 => n1441, A3 => n1442, A4 => n1443,
                           ZN => n1439);
   U501 : OAI221_X1 port map( B1 => n4943, B2 => n1453, C1 => n4940, C2 => 
                           n1454, A => n1455, ZN => n1440);
   U502 : OAI221_X1 port map( B1 => n4955, B2 => n1450, C1 => n4952, C2 => 
                           n1451, A => n1452, ZN => n1441);
   U503 : OAI221_X1 port map( B1 => n4967, B2 => n1447, C1 => n4964, C2 => 
                           n1448, A => n1449, ZN => n1442);
   U504 : NOR4_X1 port map( A1 => n1407, A2 => n1408, A3 => n1409, A4 => n1410,
                           ZN => n1406);
   U505 : OAI221_X1 port map( B1 => n4943, B2 => n1420, C1 => n4940, C2 => 
                           n1421, A => n1422, ZN => n1407);
   U506 : OAI221_X1 port map( B1 => n4955, B2 => n1417, C1 => n4952, C2 => 
                           n1418, A => n1419, ZN => n1408);
   U507 : OAI221_X1 port map( B1 => n4967, B2 => n1414, C1 => n4964, C2 => 
                           n1415, A => n1416, ZN => n1409);
   U508 : NOR4_X1 port map( A1 => n1374, A2 => n1375, A3 => n1376, A4 => n1377,
                           ZN => n1373);
   U509 : OAI221_X1 port map( B1 => n4943, B2 => n1387, C1 => n4940, C2 => 
                           n1388, A => n1389, ZN => n1374);
   U510 : OAI221_X1 port map( B1 => n4955, B2 => n1384, C1 => n4952, C2 => 
                           n1385, A => n1386, ZN => n1375);
   U511 : OAI221_X1 port map( B1 => n4967, B2 => n1381, C1 => n4964, C2 => 
                           n1382, A => n1383, ZN => n1376);
   U512 : NOR4_X1 port map( A1 => n1341, A2 => n1342, A3 => n1343, A4 => n1344,
                           ZN => n1340);
   U513 : OAI221_X1 port map( B1 => n4943, B2 => n1354, C1 => n4940, C2 => 
                           n1355, A => n1356, ZN => n1341);
   U514 : OAI221_X1 port map( B1 => n4955, B2 => n1351, C1 => n4952, C2 => 
                           n1352, A => n1353, ZN => n1342);
   U515 : OAI221_X1 port map( B1 => n4967, B2 => n1348, C1 => n4964, C2 => 
                           n1349, A => n1350, ZN => n1343);
   U516 : NOR4_X1 port map( A1 => n1308, A2 => n1309, A3 => n1310, A4 => n1311,
                           ZN => n1307);
   U517 : OAI221_X1 port map( B1 => n4943, B2 => n1321, C1 => n4940, C2 => 
                           n1322, A => n1323, ZN => n1308);
   U518 : OAI221_X1 port map( B1 => n4955, B2 => n1318, C1 => n4952, C2 => 
                           n1319, A => n1320, ZN => n1309);
   U519 : OAI221_X1 port map( B1 => n4967, B2 => n1315, C1 => n4964, C2 => 
                           n1316, A => n1317, ZN => n1310);
   U520 : NOR4_X1 port map( A1 => n1275, A2 => n1276, A3 => n1277, A4 => n1278,
                           ZN => n1274);
   U521 : OAI221_X1 port map( B1 => n4943, B2 => n1288, C1 => n4940, C2 => 
                           n1289, A => n1290, ZN => n1275);
   U522 : OAI221_X1 port map( B1 => n4955, B2 => n1285, C1 => n4952, C2 => 
                           n1286, A => n1287, ZN => n1276);
   U523 : OAI221_X1 port map( B1 => n4967, B2 => n1282, C1 => n4964, C2 => 
                           n1283, A => n1284, ZN => n1277);
   U524 : NOR4_X1 port map( A1 => n1242, A2 => n1243, A3 => n1244, A4 => n1245,
                           ZN => n1241);
   U525 : OAI221_X1 port map( B1 => n4943, B2 => n1255, C1 => n4940, C2 => 
                           n1256, A => n1257, ZN => n1242);
   U526 : OAI221_X1 port map( B1 => n4955, B2 => n1252, C1 => n4952, C2 => 
                           n1253, A => n1254, ZN => n1243);
   U527 : OAI221_X1 port map( B1 => n4967, B2 => n1249, C1 => n4964, C2 => 
                           n1250, A => n1251, ZN => n1244);
   U528 : NOR4_X1 port map( A1 => n1209, A2 => n1210, A3 => n1211, A4 => n1212,
                           ZN => n1208);
   U529 : OAI221_X1 port map( B1 => n4944, B2 => n1222, C1 => n4941, C2 => 
                           n1223, A => n1224, ZN => n1209);
   U530 : OAI221_X1 port map( B1 => n4956, B2 => n1219, C1 => n4953, C2 => 
                           n1220, A => n1221, ZN => n1210);
   U531 : OAI221_X1 port map( B1 => n4968, B2 => n1216, C1 => n4965, C2 => 
                           n1217, A => n1218, ZN => n1211);
   U532 : NOR4_X1 port map( A1 => n1176, A2 => n1177, A3 => n1178, A4 => n1179,
                           ZN => n1175);
   U533 : OAI221_X1 port map( B1 => n4944, B2 => n1189, C1 => n4941, C2 => 
                           n1190, A => n1191, ZN => n1176);
   U534 : OAI221_X1 port map( B1 => n4956, B2 => n1186, C1 => n4953, C2 => 
                           n1187, A => n1188, ZN => n1177);
   U535 : OAI221_X1 port map( B1 => n4968, B2 => n1183, C1 => n4965, C2 => 
                           n1184, A => n1185, ZN => n1178);
   U536 : NOR4_X1 port map( A1 => n1143, A2 => n1144, A3 => n1145, A4 => n1146,
                           ZN => n1142);
   U537 : OAI221_X1 port map( B1 => n4944, B2 => n1156, C1 => n4941, C2 => 
                           n1157, A => n1158, ZN => n1143);
   U538 : OAI221_X1 port map( B1 => n4956, B2 => n1153, C1 => n4953, C2 => 
                           n1154, A => n1155, ZN => n1144);
   U539 : OAI221_X1 port map( B1 => n4968, B2 => n1150, C1 => n4965, C2 => 
                           n1151, A => n1152, ZN => n1145);
   U540 : NOR4_X1 port map( A1 => n1110, A2 => n1111, A3 => n1112, A4 => n1113,
                           ZN => n1109);
   U541 : OAI221_X1 port map( B1 => n4944, B2 => n1123, C1 => n4941, C2 => 
                           n1124, A => n1125, ZN => n1110);
   U542 : OAI221_X1 port map( B1 => n4956, B2 => n1120, C1 => n4953, C2 => 
                           n1121, A => n1122, ZN => n1111);
   U543 : OAI221_X1 port map( B1 => n4968, B2 => n1117, C1 => n4965, C2 => 
                           n1118, A => n1119, ZN => n1112);
   U544 : OAI21_X1 port map( B1 => n540, B2 => n541, A => n5178, ZN => n2952);
   U545 : OAI21_X1 port map( B1 => n530, B2 => n537, A => n5179, ZN => n2955);
   U546 : OAI21_X1 port map( B1 => n530, B2 => n536, A => n5179, ZN => n2958);
   U547 : OAI21_X1 port map( B1 => n530, B2 => n535, A => n5179, ZN => n2961);
   U548 : OAI21_X1 port map( B1 => n530, B2 => n534, A => n5179, ZN => n2964);
   U549 : OAI21_X1 port map( B1 => n530, B2 => n533, A => n5179, ZN => n2967);
   U550 : OAI21_X1 port map( B1 => n530, B2 => n532, A => n5179, ZN => n2970);
   U551 : OAI21_X1 port map( B1 => n530, B2 => n531, A => n5179, ZN => n2973);
   U552 : OAI22_X1 port map( A1 => n4906, A2 => n837, B1 => n4903, B2 => n838, 
                           ZN => n836);
   U553 : OAI22_X1 port map( A1 => n4894, A2 => n840, B1 => n4891, B2 => n841, 
                           ZN => n839);
   U554 : OAI22_X1 port map( A1 => n4906, A2 => n804, B1 => n4903, B2 => n805, 
                           ZN => n803);
   U555 : OAI22_X1 port map( A1 => n4894, A2 => n807, B1 => n4891, B2 => n808, 
                           ZN => n806);
   U556 : OAI22_X1 port map( A1 => n4906, A2 => n771, B1 => n4903, B2 => n772, 
                           ZN => n770);
   U557 : OAI22_X1 port map( A1 => n4894, A2 => n774, B1 => n4891, B2 => n775, 
                           ZN => n773);
   U558 : OAI22_X1 port map( A1 => n4906, A2 => n738, B1 => n4903, B2 => n739, 
                           ZN => n737);
   U559 : OAI22_X1 port map( A1 => n4894, A2 => n741, B1 => n4891, B2 => n742, 
                           ZN => n740);
   U560 : OAI22_X1 port map( A1 => n4906, A2 => n705, B1 => n4903, B2 => n706, 
                           ZN => n704);
   U561 : OAI22_X1 port map( A1 => n4894, A2 => n708, B1 => n4891, B2 => n709, 
                           ZN => n707);
   U562 : OAI22_X1 port map( A1 => n4906, A2 => n672, B1 => n4903, B2 => n673, 
                           ZN => n671);
   U563 : OAI22_X1 port map( A1 => n4894, A2 => n675, B1 => n4891, B2 => n676, 
                           ZN => n674);
   U564 : OAI22_X1 port map( A1 => n4906, A2 => n639, B1 => n4903, B2 => n640, 
                           ZN => n638);
   U565 : OAI22_X1 port map( A1 => n4894, A2 => n642, B1 => n4891, B2 => n643, 
                           ZN => n641);
   U566 : OAI22_X1 port map( A1 => n4906, A2 => n601, B1 => n4903, B2 => n603, 
                           ZN => n599);
   U567 : OAI22_X1 port map( A1 => n4894, A2 => n608, B1 => n4891, B2 => n610, 
                           ZN => n606);
   U568 : OAI22_X1 port map( A1 => n4930, A2 => n831, B1 => n4927, B2 => n832, 
                           ZN => n830);
   U569 : OAI22_X1 port map( A1 => n4930, A2 => n798, B1 => n4927, B2 => n799, 
                           ZN => n797);
   U570 : OAI22_X1 port map( A1 => n4930, A2 => n765, B1 => n4927, B2 => n766, 
                           ZN => n764);
   U571 : OAI22_X1 port map( A1 => n4930, A2 => n732, B1 => n4927, B2 => n733, 
                           ZN => n731);
   U572 : OAI22_X1 port map( A1 => n4930, A2 => n699, B1 => n4927, B2 => n700, 
                           ZN => n698);
   U573 : OAI22_X1 port map( A1 => n4930, A2 => n666, B1 => n4927, B2 => n667, 
                           ZN => n665);
   U574 : OAI22_X1 port map( A1 => n4930, A2 => n633, B1 => n4927, B2 => n634, 
                           ZN => n632);
   U575 : OAI22_X1 port map( A1 => n4930, A2 => n587, B1 => n4927, B2 => n589, 
                           ZN => n585);
   U576 : OAI22_X1 port map( A1 => n837, A2 => n4813, B1 => n838, B2 => n4810, 
                           ZN => n1880);
   U577 : OAI22_X1 port map( A1 => n840, A2 => n4801, B1 => n841, B2 => n4798, 
                           ZN => n1881);
   U578 : OAI22_X1 port map( A1 => n804, A2 => n4813, B1 => n805, B2 => n4810, 
                           ZN => n1863);
   U579 : OAI22_X1 port map( A1 => n807, A2 => n4801, B1 => n808, B2 => n4798, 
                           ZN => n1864);
   U580 : OAI22_X1 port map( A1 => n771, A2 => n4813, B1 => n772, B2 => n4810, 
                           ZN => n1846);
   U581 : OAI22_X1 port map( A1 => n774, A2 => n4801, B1 => n775, B2 => n4798, 
                           ZN => n1847);
   U582 : OAI22_X1 port map( A1 => n738, A2 => n4813, B1 => n739, B2 => n4810, 
                           ZN => n1765);
   U583 : OAI22_X1 port map( A1 => n741, A2 => n4801, B1 => n742, B2 => n4798, 
                           ZN => n1766);
   U584 : OAI22_X1 port map( A1 => n705, A2 => n4813, B1 => n706, B2 => n4810, 
                           ZN => n1748);
   U585 : OAI22_X1 port map( A1 => n708, A2 => n4801, B1 => n709, B2 => n4798, 
                           ZN => n1749);
   U586 : OAI22_X1 port map( A1 => n672, A2 => n4813, B1 => n673, B2 => n4810, 
                           ZN => n1731);
   U587 : OAI22_X1 port map( A1 => n675, A2 => n4801, B1 => n676, B2 => n4798, 
                           ZN => n1732);
   U588 : OAI22_X1 port map( A1 => n639, A2 => n4813, B1 => n640, B2 => n4810, 
                           ZN => n1714);
   U589 : OAI22_X1 port map( A1 => n642, A2 => n4801, B1 => n643, B2 => n4798, 
                           ZN => n1715);
   U590 : OAI22_X1 port map( A1 => n601, A2 => n4813, B1 => n603, B2 => n4810, 
                           ZN => n1691);
   U591 : OAI22_X1 port map( A1 => n608, A2 => n4801, B1 => n610, B2 => n4798, 
                           ZN => n1696);
   U592 : OAI22_X1 port map( A1 => n831, A2 => n4837, B1 => n832, B2 => n4834, 
                           ZN => n1878);
   U593 : OAI22_X1 port map( A1 => n798, A2 => n4837, B1 => n799, B2 => n4834, 
                           ZN => n1861);
   U594 : OAI22_X1 port map( A1 => n765, A2 => n4837, B1 => n766, B2 => n4834, 
                           ZN => n1844);
   U595 : OAI22_X1 port map( A1 => n732, A2 => n4837, B1 => n733, B2 => n4834, 
                           ZN => n1763);
   U596 : OAI22_X1 port map( A1 => n699, A2 => n4837, B1 => n700, B2 => n4834, 
                           ZN => n1746);
   U597 : OAI22_X1 port map( A1 => n666, A2 => n4837, B1 => n667, B2 => n4834, 
                           ZN => n1729);
   U598 : OAI22_X1 port map( A1 => n633, A2 => n4837, B1 => n634, B2 => n4834, 
                           ZN => n1712);
   U599 : OAI22_X1 port map( A1 => n587, A2 => n4837, B1 => n589, B2 => n4834, 
                           ZN => n1681);
   U600 : OAI22_X1 port map( A1 => n1101, A2 => n4812, B1 => n1102, B2 => n4809
                           , ZN => n2016);
   U601 : OAI22_X1 port map( A1 => n1104, A2 => n4800, B1 => n1105, B2 => n4797
                           , ZN => n2017);
   U602 : OAI22_X1 port map( A1 => n1068, A2 => n4812, B1 => n1069, B2 => n4809
                           , ZN => n1999);
   U603 : OAI22_X1 port map( A1 => n1071, A2 => n4800, B1 => n1072, B2 => n4797
                           , ZN => n2000);
   U604 : OAI22_X1 port map( A1 => n1035, A2 => n4812, B1 => n1036, B2 => n4809
                           , ZN => n1982);
   U605 : OAI22_X1 port map( A1 => n1038, A2 => n4800, B1 => n1039, B2 => n4797
                           , ZN => n1983);
   U606 : OAI22_X1 port map( A1 => n1002, A2 => n4812, B1 => n1003, B2 => n4809
                           , ZN => n1965);
   U607 : OAI22_X1 port map( A1 => n1005, A2 => n4800, B1 => n1006, B2 => n4797
                           , ZN => n1966);
   U608 : OAI22_X1 port map( A1 => n969, A2 => n4812, B1 => n970, B2 => n4809, 
                           ZN => n1948);
   U609 : OAI22_X1 port map( A1 => n972, A2 => n4800, B1 => n973, B2 => n4797, 
                           ZN => n1949);
   U610 : OAI22_X1 port map( A1 => n936, A2 => n4812, B1 => n937, B2 => n4809, 
                           ZN => n1931);
   U611 : OAI22_X1 port map( A1 => n939, A2 => n4800, B1 => n940, B2 => n4797, 
                           ZN => n1932);
   U612 : OAI22_X1 port map( A1 => n903, A2 => n4812, B1 => n904, B2 => n4809, 
                           ZN => n1914);
   U613 : OAI22_X1 port map( A1 => n906, A2 => n4800, B1 => n907, B2 => n4797, 
                           ZN => n1915);
   U614 : OAI22_X1 port map( A1 => n870, A2 => n4812, B1 => n871, B2 => n4809, 
                           ZN => n1897);
   U615 : OAI22_X1 port map( A1 => n873, A2 => n4800, B1 => n874, B2 => n4797, 
                           ZN => n1898);
   U616 : OAI22_X1 port map( A1 => n4905, A2 => n1101, B1 => n4902, B2 => n1102
                           , ZN => n1100);
   U617 : OAI22_X1 port map( A1 => n4893, A2 => n1104, B1 => n4890, B2 => n1105
                           , ZN => n1103);
   U618 : OAI22_X1 port map( A1 => n4905, A2 => n1068, B1 => n4902, B2 => n1069
                           , ZN => n1067);
   U619 : OAI22_X1 port map( A1 => n4893, A2 => n1071, B1 => n4890, B2 => n1072
                           , ZN => n1070);
   U620 : OAI22_X1 port map( A1 => n4905, A2 => n1035, B1 => n4902, B2 => n1036
                           , ZN => n1034);
   U621 : OAI22_X1 port map( A1 => n4893, A2 => n1038, B1 => n4890, B2 => n1039
                           , ZN => n1037);
   U622 : OAI22_X1 port map( A1 => n4905, A2 => n1002, B1 => n4902, B2 => n1003
                           , ZN => n1001);
   U623 : OAI22_X1 port map( A1 => n4893, A2 => n1005, B1 => n4890, B2 => n1006
                           , ZN => n1004);
   U624 : OAI22_X1 port map( A1 => n4905, A2 => n969, B1 => n4902, B2 => n970, 
                           ZN => n968);
   U625 : OAI22_X1 port map( A1 => n4893, A2 => n972, B1 => n4890, B2 => n973, 
                           ZN => n971);
   U626 : OAI22_X1 port map( A1 => n4905, A2 => n936, B1 => n4902, B2 => n937, 
                           ZN => n935);
   U627 : OAI22_X1 port map( A1 => n4893, A2 => n939, B1 => n4890, B2 => n940, 
                           ZN => n938);
   U628 : OAI22_X1 port map( A1 => n4905, A2 => n903, B1 => n4902, B2 => n904, 
                           ZN => n902);
   U629 : OAI22_X1 port map( A1 => n4893, A2 => n906, B1 => n4890, B2 => n907, 
                           ZN => n905);
   U630 : OAI22_X1 port map( A1 => n4905, A2 => n870, B1 => n4902, B2 => n871, 
                           ZN => n869);
   U631 : OAI22_X1 port map( A1 => n4893, A2 => n873, B1 => n4890, B2 => n874, 
                           ZN => n872);
   U632 : OAI22_X1 port map( A1 => n1644, A2 => n4811, B1 => n1645, B2 => n4808
                           , ZN => n2303);
   U633 : OAI22_X1 port map( A1 => n1647, A2 => n4799, B1 => n1648, B2 => n4796
                           , ZN => n2304);
   U634 : OAI22_X1 port map( A1 => n1596, A2 => n4811, B1 => n1597, B2 => n4808
                           , ZN => n2271);
   U635 : OAI22_X1 port map( A1 => n1599, A2 => n4799, B1 => n1600, B2 => n4796
                           , ZN => n2272);
   U636 : OAI22_X1 port map( A1 => n1563, A2 => n4811, B1 => n1564, B2 => n4808
                           , ZN => n2254);
   U637 : OAI22_X1 port map( A1 => n1566, A2 => n4799, B1 => n1567, B2 => n4796
                           , ZN => n2255);
   U638 : OAI22_X1 port map( A1 => n1530, A2 => n4811, B1 => n1531, B2 => n4808
                           , ZN => n2237);
   U639 : OAI22_X1 port map( A1 => n1533, A2 => n4799, B1 => n1534, B2 => n4796
                           , ZN => n2238);
   U640 : OAI22_X1 port map( A1 => n1497, A2 => n4811, B1 => n1498, B2 => n4808
                           , ZN => n2220);
   U641 : OAI22_X1 port map( A1 => n1500, A2 => n4799, B1 => n1501, B2 => n4796
                           , ZN => n2221);
   U642 : OAI22_X1 port map( A1 => n1464, A2 => n4811, B1 => n1465, B2 => n4808
                           , ZN => n2203);
   U643 : OAI22_X1 port map( A1 => n1467, A2 => n4799, B1 => n1468, B2 => n4796
                           , ZN => n2204);
   U644 : OAI22_X1 port map( A1 => n1431, A2 => n4811, B1 => n1432, B2 => n4808
                           , ZN => n2186);
   U645 : OAI22_X1 port map( A1 => n1434, A2 => n4799, B1 => n1435, B2 => n4796
                           , ZN => n2187);
   U646 : OAI22_X1 port map( A1 => n1398, A2 => n4811, B1 => n1399, B2 => n4808
                           , ZN => n2169);
   U647 : OAI22_X1 port map( A1 => n1401, A2 => n4799, B1 => n1402, B2 => n4796
                           , ZN => n2170);
   U648 : OAI22_X1 port map( A1 => n1365, A2 => n4811, B1 => n1366, B2 => n4808
                           , ZN => n2152);
   U649 : OAI22_X1 port map( A1 => n1368, A2 => n4799, B1 => n1369, B2 => n4796
                           , ZN => n2153);
   U650 : OAI22_X1 port map( A1 => n1332, A2 => n4811, B1 => n1333, B2 => n4808
                           , ZN => n2135);
   U651 : OAI22_X1 port map( A1 => n1335, A2 => n4799, B1 => n1336, B2 => n4796
                           , ZN => n2136);
   U652 : OAI22_X1 port map( A1 => n1299, A2 => n4811, B1 => n1300, B2 => n4808
                           , ZN => n2118);
   U653 : OAI22_X1 port map( A1 => n1302, A2 => n4799, B1 => n1303, B2 => n4796
                           , ZN => n2119);
   U654 : OAI22_X1 port map( A1 => n1266, A2 => n4811, B1 => n1267, B2 => n4808
                           , ZN => n2101);
   U655 : OAI22_X1 port map( A1 => n1269, A2 => n4799, B1 => n1270, B2 => n4796
                           , ZN => n2102);
   U656 : OAI22_X1 port map( A1 => n1233, A2 => n4812, B1 => n1234, B2 => n4809
                           , ZN => n2084);
   U657 : OAI22_X1 port map( A1 => n1236, A2 => n4800, B1 => n1237, B2 => n4797
                           , ZN => n2085);
   U658 : OAI22_X1 port map( A1 => n1200, A2 => n4812, B1 => n1201, B2 => n4809
                           , ZN => n2067);
   U659 : OAI22_X1 port map( A1 => n1203, A2 => n4800, B1 => n1204, B2 => n4797
                           , ZN => n2068);
   U660 : OAI22_X1 port map( A1 => n1167, A2 => n4812, B1 => n1168, B2 => n4809
                           , ZN => n2050);
   U661 : OAI22_X1 port map( A1 => n1170, A2 => n4800, B1 => n1171, B2 => n4797
                           , ZN => n2051);
   U662 : OAI22_X1 port map( A1 => n1134, A2 => n4812, B1 => n1135, B2 => n4809
                           , ZN => n2033);
   U663 : OAI22_X1 port map( A1 => n1137, A2 => n4800, B1 => n1138, B2 => n4797
                           , ZN => n2034);
   U664 : OAI22_X1 port map( A1 => n4904, A2 => n1644, B1 => n4901, B2 => n1645
                           , ZN => n1643);
   U665 : OAI22_X1 port map( A1 => n4892, A2 => n1647, B1 => n4889, B2 => n1648
                           , ZN => n1646);
   U666 : OAI22_X1 port map( A1 => n4904, A2 => n1596, B1 => n4901, B2 => n1597
                           , ZN => n1595);
   U667 : OAI22_X1 port map( A1 => n4892, A2 => n1599, B1 => n4889, B2 => n1600
                           , ZN => n1598);
   U668 : OAI22_X1 port map( A1 => n4904, A2 => n1563, B1 => n4901, B2 => n1564
                           , ZN => n1562);
   U669 : OAI22_X1 port map( A1 => n4892, A2 => n1566, B1 => n4889, B2 => n1567
                           , ZN => n1565);
   U670 : OAI22_X1 port map( A1 => n4904, A2 => n1530, B1 => n4901, B2 => n1531
                           , ZN => n1529);
   U671 : OAI22_X1 port map( A1 => n4892, A2 => n1533, B1 => n4889, B2 => n1534
                           , ZN => n1532);
   U672 : OAI22_X1 port map( A1 => n4904, A2 => n1497, B1 => n4901, B2 => n1498
                           , ZN => n1496);
   U673 : OAI22_X1 port map( A1 => n4892, A2 => n1500, B1 => n4889, B2 => n1501
                           , ZN => n1499);
   U674 : OAI22_X1 port map( A1 => n4904, A2 => n1464, B1 => n4901, B2 => n1465
                           , ZN => n1463);
   U675 : OAI22_X1 port map( A1 => n4892, A2 => n1467, B1 => n4889, B2 => n1468
                           , ZN => n1466);
   U676 : OAI22_X1 port map( A1 => n4904, A2 => n1431, B1 => n4901, B2 => n1432
                           , ZN => n1430);
   U677 : OAI22_X1 port map( A1 => n4892, A2 => n1434, B1 => n4889, B2 => n1435
                           , ZN => n1433);
   U678 : OAI22_X1 port map( A1 => n4904, A2 => n1398, B1 => n4901, B2 => n1399
                           , ZN => n1397);
   U679 : OAI22_X1 port map( A1 => n4892, A2 => n1401, B1 => n4889, B2 => n1402
                           , ZN => n1400);
   U680 : OAI22_X1 port map( A1 => n4904, A2 => n1365, B1 => n4901, B2 => n1366
                           , ZN => n1364);
   U681 : OAI22_X1 port map( A1 => n4892, A2 => n1368, B1 => n4889, B2 => n1369
                           , ZN => n1367);
   U682 : OAI22_X1 port map( A1 => n4904, A2 => n1332, B1 => n4901, B2 => n1333
                           , ZN => n1331);
   U683 : OAI22_X1 port map( A1 => n4892, A2 => n1335, B1 => n4889, B2 => n1336
                           , ZN => n1334);
   U684 : OAI22_X1 port map( A1 => n4904, A2 => n1299, B1 => n4901, B2 => n1300
                           , ZN => n1298);
   U685 : OAI22_X1 port map( A1 => n4892, A2 => n1302, B1 => n4889, B2 => n1303
                           , ZN => n1301);
   U686 : OAI22_X1 port map( A1 => n4904, A2 => n1266, B1 => n4901, B2 => n1267
                           , ZN => n1265);
   U687 : OAI22_X1 port map( A1 => n4892, A2 => n1269, B1 => n4889, B2 => n1270
                           , ZN => n1268);
   U688 : OAI22_X1 port map( A1 => n4905, A2 => n1233, B1 => n4902, B2 => n1234
                           , ZN => n1232);
   U689 : OAI22_X1 port map( A1 => n4893, A2 => n1236, B1 => n4890, B2 => n1237
                           , ZN => n1235);
   U690 : OAI22_X1 port map( A1 => n4905, A2 => n1200, B1 => n4902, B2 => n1201
                           , ZN => n1199);
   U691 : OAI22_X1 port map( A1 => n4893, A2 => n1203, B1 => n4890, B2 => n1204
                           , ZN => n1202);
   U692 : OAI22_X1 port map( A1 => n4905, A2 => n1167, B1 => n4902, B2 => n1168
                           , ZN => n1166);
   U693 : OAI22_X1 port map( A1 => n4893, A2 => n1170, B1 => n4890, B2 => n1171
                           , ZN => n1169);
   U694 : OAI22_X1 port map( A1 => n4905, A2 => n1134, B1 => n4902, B2 => n1135
                           , ZN => n1133);
   U695 : OAI22_X1 port map( A1 => n4893, A2 => n1137, B1 => n4890, B2 => n1138
                           , ZN => n1136);
   U696 : OAI21_X1 port map( B1 => n537, B2 => n543, A => n5177, ZN => n2883);
   U697 : OAI21_X1 port map( B1 => n536, B2 => n543, A => n5177, ZN => n2886);
   U698 : OAI21_X1 port map( B1 => n535, B2 => n543, A => n5177, ZN => n2889);
   U699 : OAI21_X1 port map( B1 => n534, B2 => n543, A => n5177, ZN => n2892);
   U700 : OAI21_X1 port map( B1 => n533, B2 => n543, A => n5177, ZN => n2895);
   U701 : OAI21_X1 port map( B1 => n532, B2 => n543, A => n5177, ZN => n2898);
   U702 : OAI21_X1 port map( B1 => n531, B2 => n543, A => n5177, ZN => n2901);
   U703 : OAI21_X1 port map( B1 => n541, B2 => n543, A => n5177, ZN => n2904);
   U704 : OAI21_X1 port map( B1 => n537, B2 => n542, A => n5177, ZN => n2907);
   U705 : OAI21_X1 port map( B1 => n536, B2 => n542, A => n5177, ZN => n2910);
   U706 : OAI21_X1 port map( B1 => n535, B2 => n542, A => n5177, ZN => n2913);
   U707 : OAI21_X1 port map( B1 => n534, B2 => n542, A => n5177, ZN => n2916);
   U708 : OAI21_X1 port map( B1 => n533, B2 => n542, A => n5178, ZN => n2919);
   U709 : OAI21_X1 port map( B1 => n532, B2 => n542, A => n5178, ZN => n2922);
   U710 : OAI21_X1 port map( B1 => n531, B2 => n542, A => n5178, ZN => n2925);
   U711 : OAI21_X1 port map( B1 => n541, B2 => n542, A => n5178, ZN => n2928);
   U712 : OAI22_X1 port map( A1 => n1095, A2 => n4836, B1 => n1096, B2 => n4833
                           , ZN => n2014);
   U713 : OAI22_X1 port map( A1 => n1062, A2 => n4836, B1 => n1063, B2 => n4833
                           , ZN => n1997);
   U714 : OAI22_X1 port map( A1 => n1029, A2 => n4836, B1 => n1030, B2 => n4833
                           , ZN => n1980);
   U715 : OAI22_X1 port map( A1 => n996, A2 => n4836, B1 => n997, B2 => n4833, 
                           ZN => n1963);
   U716 : OAI22_X1 port map( A1 => n963, A2 => n4836, B1 => n964, B2 => n4833, 
                           ZN => n1946);
   U717 : OAI22_X1 port map( A1 => n930, A2 => n4836, B1 => n931, B2 => n4833, 
                           ZN => n1929);
   U718 : OAI22_X1 port map( A1 => n897, A2 => n4836, B1 => n898, B2 => n4833, 
                           ZN => n1912);
   U719 : OAI22_X1 port map( A1 => n864, A2 => n4836, B1 => n865, B2 => n4833, 
                           ZN => n1895);
   U720 : OAI22_X1 port map( A1 => n4929, A2 => n1095, B1 => n4926, B2 => n1096
                           , ZN => n1094);
   U721 : OAI22_X1 port map( A1 => n4929, A2 => n1062, B1 => n4926, B2 => n1063
                           , ZN => n1061);
   U722 : OAI22_X1 port map( A1 => n4929, A2 => n1029, B1 => n4926, B2 => n1030
                           , ZN => n1028);
   U723 : OAI22_X1 port map( A1 => n4929, A2 => n996, B1 => n4926, B2 => n997, 
                           ZN => n995);
   U724 : OAI22_X1 port map( A1 => n4929, A2 => n963, B1 => n4926, B2 => n964, 
                           ZN => n962);
   U725 : OAI22_X1 port map( A1 => n4929, A2 => n930, B1 => n4926, B2 => n931, 
                           ZN => n929);
   U726 : OAI22_X1 port map( A1 => n4929, A2 => n897, B1 => n4926, B2 => n898, 
                           ZN => n896);
   U727 : OAI22_X1 port map( A1 => n4929, A2 => n864, B1 => n4926, B2 => n865, 
                           ZN => n863);
   U728 : OAI22_X1 port map( A1 => n1635, A2 => n4835, B1 => n1636, B2 => n4832
                           , ZN => n2298);
   U729 : OAI22_X1 port map( A1 => n1590, A2 => n4835, B1 => n1591, B2 => n4832
                           , ZN => n2269);
   U730 : OAI22_X1 port map( A1 => n1557, A2 => n4835, B1 => n1558, B2 => n4832
                           , ZN => n2252);
   U731 : OAI22_X1 port map( A1 => n1524, A2 => n4835, B1 => n1525, B2 => n4832
                           , ZN => n2235);
   U732 : OAI22_X1 port map( A1 => n1491, A2 => n4835, B1 => n1492, B2 => n4832
                           , ZN => n2218);
   U733 : OAI22_X1 port map( A1 => n1458, A2 => n4835, B1 => n1459, B2 => n4832
                           , ZN => n2201);
   U734 : OAI22_X1 port map( A1 => n1425, A2 => n4835, B1 => n1426, B2 => n4832
                           , ZN => n2184);
   U735 : OAI22_X1 port map( A1 => n1392, A2 => n4835, B1 => n1393, B2 => n4832
                           , ZN => n2167);
   U736 : OAI22_X1 port map( A1 => n1359, A2 => n4835, B1 => n1360, B2 => n4832
                           , ZN => n2150);
   U737 : OAI22_X1 port map( A1 => n1326, A2 => n4835, B1 => n1327, B2 => n4832
                           , ZN => n2133);
   U738 : OAI22_X1 port map( A1 => n1293, A2 => n4835, B1 => n1294, B2 => n4832
                           , ZN => n2116);
   U739 : OAI22_X1 port map( A1 => n1260, A2 => n4835, B1 => n1261, B2 => n4832
                           , ZN => n2099);
   U740 : OAI22_X1 port map( A1 => n1227, A2 => n4836, B1 => n1228, B2 => n4833
                           , ZN => n2082);
   U741 : OAI22_X1 port map( A1 => n1194, A2 => n4836, B1 => n1195, B2 => n4833
                           , ZN => n2065);
   U742 : OAI22_X1 port map( A1 => n1161, A2 => n4836, B1 => n1162, B2 => n4833
                           , ZN => n2048);
   U743 : OAI22_X1 port map( A1 => n1128, A2 => n4836, B1 => n1129, B2 => n4833
                           , ZN => n2031);
   U744 : OAI22_X1 port map( A1 => n4928, A2 => n1635, B1 => n4925, B2 => n1636
                           , ZN => n1634);
   U745 : OAI22_X1 port map( A1 => n4928, A2 => n1590, B1 => n4925, B2 => n1591
                           , ZN => n1589);
   U746 : OAI22_X1 port map( A1 => n4928, A2 => n1557, B1 => n4925, B2 => n1558
                           , ZN => n1556);
   U747 : OAI22_X1 port map( A1 => n4928, A2 => n1524, B1 => n4925, B2 => n1525
                           , ZN => n1523);
   U748 : OAI22_X1 port map( A1 => n4928, A2 => n1491, B1 => n4925, B2 => n1492
                           , ZN => n1490);
   U749 : OAI22_X1 port map( A1 => n4928, A2 => n1458, B1 => n4925, B2 => n1459
                           , ZN => n1457);
   U750 : OAI22_X1 port map( A1 => n4928, A2 => n1425, B1 => n4925, B2 => n1426
                           , ZN => n1424);
   U751 : OAI22_X1 port map( A1 => n4928, A2 => n1392, B1 => n4925, B2 => n1393
                           , ZN => n1391);
   U752 : OAI22_X1 port map( A1 => n4928, A2 => n1359, B1 => n4925, B2 => n1360
                           , ZN => n1358);
   U753 : OAI22_X1 port map( A1 => n4928, A2 => n1326, B1 => n4925, B2 => n1327
                           , ZN => n1325);
   U754 : OAI22_X1 port map( A1 => n4928, A2 => n1293, B1 => n4925, B2 => n1294
                           , ZN => n1292);
   U755 : OAI22_X1 port map( A1 => n4928, A2 => n1260, B1 => n4925, B2 => n1261
                           , ZN => n1259);
   U756 : OAI22_X1 port map( A1 => n4929, A2 => n1227, B1 => n4926, B2 => n1228
                           , ZN => n1226);
   U757 : OAI22_X1 port map( A1 => n4929, A2 => n1194, B1 => n4926, B2 => n1195
                           , ZN => n1193);
   U758 : OAI22_X1 port map( A1 => n4929, A2 => n1161, B1 => n4926, B2 => n1162
                           , ZN => n1160);
   U759 : OAI22_X1 port map( A1 => n4929, A2 => n1128, B1 => n4926, B2 => n1129
                           , ZN => n1127);
   U760 : OAI21_X1 port map( B1 => n537, B2 => n540, A => n5178, ZN => n2931);
   U761 : OAI21_X1 port map( B1 => n536, B2 => n540, A => n5178, ZN => n2934);
   U762 : OAI21_X1 port map( B1 => n535, B2 => n540, A => n5178, ZN => n2937);
   U763 : OAI21_X1 port map( B1 => n534, B2 => n540, A => n5178, ZN => n2940);
   U764 : OAI21_X1 port map( B1 => n533, B2 => n540, A => n5178, ZN => n2943);
   U765 : OAI21_X1 port map( B1 => n532, B2 => n540, A => n5178, ZN => n2946);
   U766 : OAI21_X1 port map( B1 => n531, B2 => n540, A => n5178, ZN => n2949);
   U767 : BUF_X1 port map( A => n5182, Z => n5179);
   U768 : BUF_X1 port map( A => n5182, Z => n5177);
   U769 : BUF_X1 port map( A => n5182, Z => n5178);
   U770 : BUF_X1 port map( A => n5182, Z => n5180);
   U771 : BUF_X1 port map( A => n3072, Z => n4985);
   U772 : BUF_X1 port map( A => n3075, Z => n4982);
   U773 : BUF_X1 port map( A => n3072, Z => n4986);
   U774 : BUF_X1 port map( A => n3075, Z => n4983);
   U775 : BUF_X1 port map( A => n3072, Z => n4987);
   U776 : BUF_X1 port map( A => n3075, Z => n4984);
   U777 : NAND2_X1 port map( A1 => n2282, A2 => n2295, ZN => n1693);
   U778 : NAND2_X1 port map( A1 => n2282, A2 => n2290, ZN => n1698);
   U779 : NAND2_X1 port map( A1 => n2282, A2 => n2292, ZN => n1685);
   U780 : NAND2_X1 port map( A1 => n2282, A2 => n2284, ZN => n1684);
   U781 : NAND2_X1 port map( A1 => n2282, A2 => n2294, ZN => n1683);
   U782 : NAND2_X1 port map( A1 => n1612, A2 => n1629, ZN => n602);
   U783 : NAND2_X1 port map( A1 => n1612, A2 => n1622, ZN => n609);
   U784 : NAND2_X1 port map( A1 => n1612, A2 => n1614, ZN => n590);
   U785 : NAND2_X1 port map( A1 => n1612, A2 => n1624, ZN => n592);
   U786 : NAND2_X1 port map( A1 => n1612, A2 => n1628, ZN => n588);
   U787 : NAND2_X1 port map( A1 => n2294, A2 => n2286, ZN => n1675);
   U788 : NAND2_X1 port map( A1 => n1628, A2 => n1616, ZN => n578);
   U789 : NAND2_X1 port map( A1 => n1624, A2 => n1615, ZN => n562);
   U790 : NAND2_X1 port map( A1 => n1624, A2 => n1616, ZN => n571);
   U791 : NAND2_X1 port map( A1 => n2292, A2 => n2285, ZN => n1664);
   U792 : NAND2_X1 port map( A1 => n2292, A2 => n2286, ZN => n1670);
   U793 : NAND2_X1 port map( A1 => n2287, A2 => n2295, ZN => n1692);
   U794 : NAND2_X1 port map( A1 => n2287, A2 => n2294, ZN => n1697);
   U795 : NAND2_X1 port map( A1 => n2287, A2 => n2283, ZN => n1682);
   U796 : NAND2_X1 port map( A1 => n1617, A2 => n1629, ZN => n600);
   U797 : NAND2_X1 port map( A1 => n1617, A2 => n1628, ZN => n607);
   U798 : NAND2_X1 port map( A1 => n1617, A2 => n1613, ZN => n586);
   U799 : NAND2_X1 port map( A1 => n1613, A2 => n1616, ZN => n576);
   U800 : NAND2_X1 port map( A1 => n2283, A2 => n2286, ZN => n1674);
   U801 : NAND2_X1 port map( A1 => n1614, A2 => n1616, ZN => n557);
   U802 : NAND2_X1 port map( A1 => n2284, A2 => n2286, ZN => n1660);
   U803 : NAND2_X1 port map( A1 => n2285, A2 => n2295, ZN => n1669);
   U804 : NAND2_X1 port map( A1 => n1615, A2 => n1629, ZN => n569);
   U805 : NAND2_X1 port map( A1 => n1623, A2 => n1616, ZN => n564);
   U806 : NAND2_X1 port map( A1 => n2291, A2 => n2286, ZN => n1665);
   U807 : AND2_X1 port map( A1 => n2282, A2 => n2283, ZN => n1663);
   U808 : AND2_X1 port map( A1 => n1612, A2 => n1613, ZN => n561);
   U809 : AND2_X1 port map( A1 => n2282, A2 => n2288, ZN => n1689);
   U810 : AND2_X1 port map( A1 => n2282, A2 => n2291, ZN => n1695);
   U811 : AND2_X1 port map( A1 => n1612, A2 => n1618, ZN => n597);
   U812 : AND2_X1 port map( A1 => n1612, A2 => n1623, ZN => n605);
   U813 : AND2_X1 port map( A1 => n2287, A2 => n2290, ZN => n1668);
   U814 : AND2_X1 port map( A1 => n2287, A2 => n2291, ZN => n1687);
   U815 : AND2_X1 port map( A1 => n1617, A2 => n1622, ZN => n568);
   U816 : AND2_X1 port map( A1 => n1617, A2 => n1623, ZN => n595);
   U817 : AND2_X1 port map( A1 => n2287, A2 => n2292, ZN => n1690);
   U818 : AND2_X1 port map( A1 => n1617, A2 => n1624, ZN => n598);
   U819 : AND2_X1 port map( A1 => n2284, A2 => n2285, ZN => n1662);
   U820 : AND2_X1 port map( A1 => n1614, A2 => n1615, ZN => n560);
   U821 : AND2_X1 port map( A1 => n2284, A2 => n2287, ZN => n1679);
   U822 : AND2_X1 port map( A1 => n1614, A2 => n1617, ZN => n583);
   U823 : AND2_X1 port map( A1 => n2285, A2 => n2283, ZN => n1672);
   U824 : AND2_X1 port map( A1 => n2285, A2 => n2294, ZN => n1673);
   U825 : AND2_X1 port map( A1 => n2285, A2 => n2290, ZN => n1688);
   U826 : AND2_X1 port map( A1 => n1615, A2 => n1613, ZN => n574);
   U827 : AND2_X1 port map( A1 => n1615, A2 => n1628, ZN => n575);
   U828 : AND2_X1 port map( A1 => n1615, A2 => n1622, ZN => n596);
   U829 : AND2_X1 port map( A1 => n2285, A2 => n2288, ZN => n1694);
   U830 : AND2_X1 port map( A1 => n1615, A2 => n1618, ZN => n604);
   U831 : AND2_X1 port map( A1 => n2290, A2 => n2286, ZN => n1677);
   U832 : AND2_X1 port map( A1 => n1622, A2 => n1616, ZN => n581);
   U833 : AND2_X1 port map( A1 => n2288, A2 => n2286, ZN => n1678);
   U834 : AND2_X1 port map( A1 => n1618, A2 => n1616, ZN => n582);
   U835 : AND2_X1 port map( A1 => n2291, A2 => n2285, ZN => n1667);
   U836 : AND2_X1 port map( A1 => n1623, A2 => n1615, ZN => n567);
   U837 : BUF_X1 port map( A => n2976, Z => n5081);
   U838 : BUF_X1 port map( A => n2979, Z => n5078);
   U839 : BUF_X1 port map( A => n2982, Z => n5075);
   U840 : BUF_X1 port map( A => n2985, Z => n5072);
   U841 : BUF_X1 port map( A => n2988, Z => n5069);
   U842 : BUF_X1 port map( A => n2991, Z => n5066);
   U843 : BUF_X1 port map( A => n2994, Z => n5063);
   U844 : BUF_X1 port map( A => n2997, Z => n5060);
   U845 : BUF_X1 port map( A => n3000, Z => n5057);
   U846 : BUF_X1 port map( A => n3003, Z => n5054);
   U847 : BUF_X1 port map( A => n3006, Z => n5051);
   U848 : BUF_X1 port map( A => n3009, Z => n5048);
   U849 : BUF_X1 port map( A => n3012, Z => n5045);
   U850 : BUF_X1 port map( A => n3015, Z => n5042);
   U851 : BUF_X1 port map( A => n3018, Z => n5039);
   U852 : BUF_X1 port map( A => n3021, Z => n5036);
   U853 : BUF_X1 port map( A => n3024, Z => n5033);
   U854 : BUF_X1 port map( A => n3027, Z => n5030);
   U855 : BUF_X1 port map( A => n3030, Z => n5027);
   U856 : BUF_X1 port map( A => n3033, Z => n5024);
   U857 : BUF_X1 port map( A => n3036, Z => n5021);
   U858 : BUF_X1 port map( A => n3039, Z => n5018);
   U859 : BUF_X1 port map( A => n3042, Z => n5015);
   U860 : BUF_X1 port map( A => n3045, Z => n5012);
   U861 : BUF_X1 port map( A => n3048, Z => n5009);
   U862 : BUF_X1 port map( A => n3051, Z => n5006);
   U863 : BUF_X1 port map( A => n2976, Z => n5082);
   U864 : BUF_X1 port map( A => n2979, Z => n5079);
   U865 : BUF_X1 port map( A => n2982, Z => n5076);
   U866 : BUF_X1 port map( A => n2985, Z => n5073);
   U867 : BUF_X1 port map( A => n2988, Z => n5070);
   U868 : BUF_X1 port map( A => n2991, Z => n5067);
   U869 : BUF_X1 port map( A => n2994, Z => n5064);
   U870 : BUF_X1 port map( A => n2997, Z => n5061);
   U871 : BUF_X1 port map( A => n3000, Z => n5058);
   U872 : BUF_X1 port map( A => n3003, Z => n5055);
   U873 : BUF_X1 port map( A => n3006, Z => n5052);
   U874 : BUF_X1 port map( A => n3009, Z => n5049);
   U875 : BUF_X1 port map( A => n3012, Z => n5046);
   U876 : BUF_X1 port map( A => n3015, Z => n5043);
   U877 : BUF_X1 port map( A => n3018, Z => n5040);
   U878 : BUF_X1 port map( A => n3021, Z => n5037);
   U879 : BUF_X1 port map( A => n3024, Z => n5034);
   U880 : BUF_X1 port map( A => n3027, Z => n5031);
   U881 : BUF_X1 port map( A => n3030, Z => n5028);
   U882 : BUF_X1 port map( A => n3033, Z => n5025);
   U883 : BUF_X1 port map( A => n3036, Z => n5022);
   U884 : BUF_X1 port map( A => n3039, Z => n5019);
   U885 : BUF_X1 port map( A => n3042, Z => n5016);
   U886 : BUF_X1 port map( A => n3045, Z => n5013);
   U887 : BUF_X1 port map( A => n3048, Z => n5010);
   U888 : BUF_X1 port map( A => n3051, Z => n5007);
   U889 : BUF_X1 port map( A => n3054, Z => n5003);
   U890 : BUF_X1 port map( A => n3057, Z => n5000);
   U891 : BUF_X1 port map( A => n3060, Z => n4997);
   U892 : BUF_X1 port map( A => n3063, Z => n4994);
   U893 : BUF_X1 port map( A => n3066, Z => n4991);
   U894 : BUF_X1 port map( A => n3069, Z => n4988);
   U895 : BUF_X1 port map( A => n3054, Z => n5004);
   U896 : BUF_X1 port map( A => n3057, Z => n5001);
   U897 : BUF_X1 port map( A => n3060, Z => n4998);
   U898 : BUF_X1 port map( A => n3063, Z => n4995);
   U899 : BUF_X1 port map( A => n3066, Z => n4992);
   U900 : BUF_X1 port map( A => n3069, Z => n4989);
   U901 : BUF_X1 port map( A => n5182, Z => n5181);
   U902 : BUF_X1 port map( A => n2976, Z => n5083);
   U903 : BUF_X1 port map( A => n2979, Z => n5080);
   U904 : BUF_X1 port map( A => n2982, Z => n5077);
   U905 : BUF_X1 port map( A => n2985, Z => n5074);
   U906 : BUF_X1 port map( A => n2988, Z => n5071);
   U907 : BUF_X1 port map( A => n2991, Z => n5068);
   U908 : BUF_X1 port map( A => n2994, Z => n5065);
   U909 : BUF_X1 port map( A => n2997, Z => n5062);
   U910 : BUF_X1 port map( A => n3000, Z => n5059);
   U911 : BUF_X1 port map( A => n3003, Z => n5056);
   U912 : BUF_X1 port map( A => n3006, Z => n5053);
   U913 : BUF_X1 port map( A => n3009, Z => n5050);
   U914 : BUF_X1 port map( A => n3012, Z => n5047);
   U915 : BUF_X1 port map( A => n3015, Z => n5044);
   U916 : BUF_X1 port map( A => n3018, Z => n5041);
   U917 : BUF_X1 port map( A => n3021, Z => n5038);
   U918 : BUF_X1 port map( A => n3024, Z => n5035);
   U919 : BUF_X1 port map( A => n3027, Z => n5032);
   U920 : BUF_X1 port map( A => n3030, Z => n5029);
   U921 : BUF_X1 port map( A => n3033, Z => n5026);
   U922 : BUF_X1 port map( A => n3036, Z => n5023);
   U923 : BUF_X1 port map( A => n3039, Z => n5020);
   U924 : BUF_X1 port map( A => n3042, Z => n5017);
   U925 : BUF_X1 port map( A => n3045, Z => n5014);
   U926 : BUF_X1 port map( A => n3048, Z => n5011);
   U927 : BUF_X1 port map( A => n3051, Z => n5008);
   U928 : BUF_X1 port map( A => n3054, Z => n5005);
   U929 : BUF_X1 port map( A => n3057, Z => n5002);
   U930 : BUF_X1 port map( A => n3060, Z => n4999);
   U931 : BUF_X1 port map( A => n3063, Z => n4996);
   U932 : BUF_X1 port map( A => n3066, Z => n4993);
   U933 : BUF_X1 port map( A => n3069, Z => n4990);
   U934 : NOR2_X1 port map( A1 => n2305, A2 => address_port_b(2), ZN => n2282);
   U935 : NOR2_X1 port map( A1 => n1649, A2 => address_port_a(2), ZN => n1612);
   U936 : NOR2_X1 port map( A1 => address_port_b(1), A2 => address_port_b(2), 
                           ZN => n2286);
   U937 : NOR2_X1 port map( A1 => address_port_a(1), A2 => address_port_a(2), 
                           ZN => n1616);
   U938 : NOR3_X1 port map( A1 => n1637, A2 => address_port_a(3), A3 => n1642, 
                           ZN => n1628);
   U939 : NOR3_X1 port map( A1 => n2299, A2 => address_port_b(3), A3 => n2302, 
                           ZN => n2294);
   U940 : NOR3_X1 port map( A1 => address_port_a(3), A2 => address_port_a(4), 
                           A3 => n1642, ZN => n1624);
   U941 : NOR3_X1 port map( A1 => address_port_b(3), A2 => address_port_b(4), 
                           A3 => n2302, ZN => n2292);
   U942 : NOR3_X1 port map( A1 => address_port_a(0), A2 => address_port_a(3), 
                           A3 => n1637, ZN => n1613);
   U943 : NOR3_X1 port map( A1 => address_port_b(0), A2 => address_port_b(3), 
                           A3 => n2299, ZN => n2283);
   U944 : NOR3_X1 port map( A1 => address_port_a(3), A2 => address_port_a(4), 
                           A3 => address_port_a(0), ZN => n1629);
   U945 : NOR3_X1 port map( A1 => address_port_b(3), A2 => address_port_b(4), 
                           A3 => address_port_b(0), ZN => n2295);
   U946 : NOR3_X1 port map( A1 => n1641, A2 => address_port_a(4), A3 => n1642, 
                           ZN => n1614);
   U947 : NOR3_X1 port map( A1 => n2301, A2 => address_port_b(4), A3 => n2302, 
                           ZN => n2284);
   U948 : NOR2_X1 port map( A1 => n2306, A2 => address_port_b(1), ZN => n2285);
   U949 : NOR2_X1 port map( A1 => n1650, A2 => address_port_a(1), ZN => n1615);
   U950 : NOR3_X1 port map( A1 => n2301, A2 => address_port_b(0), A3 => n2299, 
                           ZN => n2290);
   U951 : NOR3_X1 port map( A1 => n1641, A2 => address_port_a(0), A3 => n1637, 
                           ZN => n1622);
   U952 : NOR3_X1 port map( A1 => address_port_a(0), A2 => address_port_a(4), 
                           A3 => n1641, ZN => n1623);
   U953 : NOR3_X1 port map( A1 => address_port_b(0), A2 => address_port_b(4), 
                           A3 => n2301, ZN => n2291);
   U954 : OAI221_X1 port map( B1 => n4981, B2 => n817, C1 => n4978, C2 => n818,
                           A => n819, ZN => n816);
   U955 : AOI22_X1 port map( A1 => registers_13_7_port, A2 => n4975, B1 => 
                           registers_18_7_port, B2 => n4972, ZN => n819);
   U956 : OAI221_X1 port map( B1 => n4981, B2 => n784, C1 => n4978, C2 => n785,
                           A => n786, ZN => n783);
   U957 : AOI22_X1 port map( A1 => registers_13_6_port, A2 => n4975, B1 => 
                           registers_18_6_port, B2 => n4972, ZN => n786);
   U958 : OAI221_X1 port map( B1 => n4981, B2 => n751, C1 => n4978, C2 => n752,
                           A => n753, ZN => n750);
   U959 : AOI22_X1 port map( A1 => registers_13_5_port, A2 => n4975, B1 => 
                           registers_18_5_port, B2 => n4972, ZN => n753);
   U960 : OAI221_X1 port map( B1 => n4981, B2 => n718, C1 => n4978, C2 => n719,
                           A => n720, ZN => n717);
   U961 : AOI22_X1 port map( A1 => registers_13_4_port, A2 => n4975, B1 => 
                           registers_18_4_port, B2 => n4972, ZN => n720);
   U962 : OAI221_X1 port map( B1 => n4981, B2 => n685, C1 => n4978, C2 => n686,
                           A => n687, ZN => n684);
   U963 : AOI22_X1 port map( A1 => registers_13_3_port, A2 => n4975, B1 => 
                           registers_18_3_port, B2 => n4972, ZN => n687);
   U964 : OAI221_X1 port map( B1 => n4981, B2 => n652, C1 => n4978, C2 => n653,
                           A => n654, ZN => n651);
   U965 : AOI22_X1 port map( A1 => registers_13_2_port, A2 => n4975, B1 => 
                           registers_18_2_port, B2 => n4972, ZN => n654);
   U966 : OAI221_X1 port map( B1 => n4981, B2 => n619, C1 => n4978, C2 => n620,
                           A => n621, ZN => n618);
   U967 : AOI22_X1 port map( A1 => registers_13_1_port, A2 => n4975, B1 => 
                           registers_18_1_port, B2 => n4972, ZN => n621);
   U968 : OAI221_X1 port map( B1 => n4981, B2 => n556, C1 => n4978, C2 => n558,
                           A => n559, ZN => n554);
   U969 : AOI22_X1 port map( A1 => registers_13_0_port, A2 => n4975, B1 => 
                           registers_18_0_port, B2 => n4972, ZN => n559);
   U970 : OAI221_X1 port map( B1 => n817, B2 => n4888, C1 => n818, C2 => n4885,
                           A => n1873, ZN => n1872);
   U971 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_7_port, B1 => 
                           n4877, B2 => registers_18_7_port, ZN => n1873);
   U972 : OAI221_X1 port map( B1 => n784, B2 => n4888, C1 => n785, C2 => n4885,
                           A => n1856, ZN => n1855);
   U973 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_6_port, B1 => 
                           n4877, B2 => registers_18_6_port, ZN => n1856);
   U974 : OAI221_X1 port map( B1 => n751, B2 => n4888, C1 => n752, C2 => n4885,
                           A => n1775, ZN => n1774);
   U975 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_5_port, B1 => 
                           n4877, B2 => registers_18_5_port, ZN => n1775);
   U976 : OAI221_X1 port map( B1 => n718, B2 => n4888, C1 => n719, C2 => n4885,
                           A => n1758, ZN => n1757);
   U977 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_4_port, B1 => 
                           n4877, B2 => registers_18_4_port, ZN => n1758);
   U978 : OAI221_X1 port map( B1 => n685, B2 => n4888, C1 => n686, C2 => n4885,
                           A => n1741, ZN => n1740);
   U979 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_3_port, B1 => 
                           n4877, B2 => registers_18_3_port, ZN => n1741);
   U980 : OAI221_X1 port map( B1 => n652, B2 => n4888, C1 => n653, C2 => n4885,
                           A => n1724, ZN => n1723);
   U981 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_2_port, B1 => 
                           n4877, B2 => registers_18_2_port, ZN => n1724);
   U982 : OAI221_X1 port map( B1 => n619, B2 => n4888, C1 => n620, C2 => n4885,
                           A => n1707, ZN => n1706);
   U983 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_1_port, B1 => 
                           n4877, B2 => registers_18_1_port, ZN => n1707);
   U984 : OAI221_X1 port map( B1 => n556, B2 => n4888, C1 => n558, C2 => n4885,
                           A => n1661, ZN => n1658);
   U985 : AOI22_X1 port map( A1 => n4882, A2 => registers_13_0_port, B1 => 
                           n4877, B2 => registers_18_0_port, ZN => n1661);
   U986 : OAI221_X1 port map( B1 => n1081, B2 => n4887, C1 => n1082, C2 => 
                           n4884, A => n2009, ZN => n2008);
   U987 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_15_port, B1 => 
                           n4878, B2 => registers_18_15_port, ZN => n2009);
   U988 : OAI221_X1 port map( B1 => n1048, B2 => n4887, C1 => n1049, C2 => 
                           n4884, A => n1992, ZN => n1991);
   U989 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_14_port, B1 => 
                           n4878, B2 => registers_18_14_port, ZN => n1992);
   U990 : OAI221_X1 port map( B1 => n1015, B2 => n4887, C1 => n1016, C2 => 
                           n4884, A => n1975, ZN => n1974);
   U991 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_13_port, B1 => 
                           n4878, B2 => registers_18_13_port, ZN => n1975);
   U992 : OAI221_X1 port map( B1 => n982, B2 => n4887, C1 => n983, C2 => n4884,
                           A => n1958, ZN => n1957);
   U993 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_12_port, B1 => 
                           n4878, B2 => registers_18_12_port, ZN => n1958);
   U994 : OAI221_X1 port map( B1 => n949, B2 => n4887, C1 => n950, C2 => n4884,
                           A => n1941, ZN => n1940);
   U995 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_11_port, B1 => 
                           n4877, B2 => registers_18_11_port, ZN => n1941);
   U996 : OAI221_X1 port map( B1 => n916, B2 => n4887, C1 => n917, C2 => n4884,
                           A => n1924, ZN => n1923);
   U997 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_10_port, B1 => 
                           n4877, B2 => registers_18_10_port, ZN => n1924);
   U998 : OAI221_X1 port map( B1 => n883, B2 => n4887, C1 => n884, C2 => n4884,
                           A => n1907, ZN => n1906);
   U999 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_9_port, B1 => 
                           n4877, B2 => registers_18_9_port, ZN => n1907);
   U1000 : OAI221_X1 port map( B1 => n850, B2 => n4887, C1 => n851, C2 => n4884
                           , A => n1890, ZN => n1889);
   U1001 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_8_port, B1 => 
                           n4877, B2 => registers_18_8_port, ZN => n1890);
   U1002 : OAI221_X1 port map( B1 => n4980, B2 => n1081, C1 => n4977, C2 => 
                           n1082, A => n1083, ZN => n1080);
   U1003 : AOI22_X1 port map( A1 => registers_13_15_port, A2 => n4974, B1 => 
                           registers_18_15_port, B2 => n4971, ZN => n1083);
   U1004 : OAI221_X1 port map( B1 => n4980, B2 => n1048, C1 => n4977, C2 => 
                           n1049, A => n1050, ZN => n1047);
   U1005 : AOI22_X1 port map( A1 => registers_13_14_port, A2 => n4974, B1 => 
                           registers_18_14_port, B2 => n4971, ZN => n1050);
   U1006 : OAI221_X1 port map( B1 => n4980, B2 => n1015, C1 => n4977, C2 => 
                           n1016, A => n1017, ZN => n1014);
   U1007 : AOI22_X1 port map( A1 => registers_13_13_port, A2 => n4974, B1 => 
                           registers_18_13_port, B2 => n4971, ZN => n1017);
   U1008 : OAI221_X1 port map( B1 => n4980, B2 => n982, C1 => n4977, C2 => n983
                           , A => n984, ZN => n981);
   U1009 : AOI22_X1 port map( A1 => registers_13_12_port, A2 => n4974, B1 => 
                           registers_18_12_port, B2 => n4971, ZN => n984);
   U1010 : OAI221_X1 port map( B1 => n4980, B2 => n949, C1 => n4977, C2 => n950
                           , A => n951, ZN => n948);
   U1011 : AOI22_X1 port map( A1 => registers_13_11_port, A2 => n4974, B1 => 
                           registers_18_11_port, B2 => n4971, ZN => n951);
   U1012 : OAI221_X1 port map( B1 => n4980, B2 => n916, C1 => n4977, C2 => n917
                           , A => n918, ZN => n915);
   U1013 : AOI22_X1 port map( A1 => registers_13_10_port, A2 => n4974, B1 => 
                           registers_18_10_port, B2 => n4971, ZN => n918);
   U1014 : OAI221_X1 port map( B1 => n4980, B2 => n883, C1 => n4977, C2 => n884
                           , A => n885, ZN => n882);
   U1015 : AOI22_X1 port map( A1 => registers_13_9_port, A2 => n4974, B1 => 
                           registers_18_9_port, B2 => n4971, ZN => n885);
   U1016 : OAI221_X1 port map( B1 => n4980, B2 => n850, C1 => n4977, C2 => n851
                           , A => n852, ZN => n849);
   U1017 : AOI22_X1 port map( A1 => registers_13_8_port, A2 => n4974, B1 => 
                           registers_18_8_port, B2 => n4971, ZN => n852);
   U1018 : OAI221_X1 port map( B1 => n1609, B2 => n4886, C1 => n1610, C2 => 
                           n4883, A => n2281, ZN => n2280);
   U1019 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_31_port, B1 => 
                           n4879, B2 => registers_18_31_port, ZN => n2281);
   U1020 : OAI221_X1 port map( B1 => n1576, B2 => n4886, C1 => n1577, C2 => 
                           n4883, A => n2264, ZN => n2263);
   U1021 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_30_port, B1 => 
                           n4879, B2 => registers_18_30_port, ZN => n2264);
   U1022 : OAI221_X1 port map( B1 => n1543, B2 => n4886, C1 => n1544, C2 => 
                           n4883, A => n2247, ZN => n2246);
   U1023 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_29_port, B1 => 
                           n4879, B2 => registers_18_29_port, ZN => n2247);
   U1024 : OAI221_X1 port map( B1 => n1510, B2 => n4886, C1 => n1511, C2 => 
                           n4883, A => n2230, ZN => n2229);
   U1025 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_28_port, B1 => 
                           n4879, B2 => registers_18_28_port, ZN => n2230);
   U1026 : OAI221_X1 port map( B1 => n1477, B2 => n4886, C1 => n1478, C2 => 
                           n4883, A => n2213, ZN => n2212);
   U1027 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_27_port, B1 => 
                           n4879, B2 => registers_18_27_port, ZN => n2213);
   U1028 : OAI221_X1 port map( B1 => n1444, B2 => n4886, C1 => n1445, C2 => 
                           n4883, A => n2196, ZN => n2195);
   U1029 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_26_port, B1 => 
                           n4879, B2 => registers_18_26_port, ZN => n2196);
   U1030 : OAI221_X1 port map( B1 => n1411, B2 => n4886, C1 => n1412, C2 => 
                           n4883, A => n2179, ZN => n2178);
   U1031 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_25_port, B1 => 
                           n4879, B2 => registers_18_25_port, ZN => n2179);
   U1032 : OAI221_X1 port map( B1 => n1378, B2 => n4886, C1 => n1379, C2 => 
                           n4883, A => n2162, ZN => n2161);
   U1033 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_24_port, B1 => 
                           n4879, B2 => registers_18_24_port, ZN => n2162);
   U1034 : OAI221_X1 port map( B1 => n1345, B2 => n4886, C1 => n1346, C2 => 
                           n4883, A => n2145, ZN => n2144);
   U1035 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_23_port, B1 => 
                           n4878, B2 => registers_18_23_port, ZN => n2145);
   U1036 : OAI221_X1 port map( B1 => n1312, B2 => n4886, C1 => n1313, C2 => 
                           n4883, A => n2128, ZN => n2127);
   U1037 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_22_port, B1 => 
                           n4878, B2 => registers_18_22_port, ZN => n2128);
   U1038 : OAI221_X1 port map( B1 => n1279, B2 => n4886, C1 => n1280, C2 => 
                           n4883, A => n2111, ZN => n2110);
   U1039 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_21_port, B1 => 
                           n4878, B2 => registers_18_21_port, ZN => n2111);
   U1040 : OAI221_X1 port map( B1 => n1246, B2 => n4886, C1 => n1247, C2 => 
                           n4883, A => n2094, ZN => n2093);
   U1041 : AOI22_X1 port map( A1 => n4880, A2 => registers_13_20_port, B1 => 
                           n4878, B2 => registers_18_20_port, ZN => n2094);
   U1042 : OAI221_X1 port map( B1 => n1213, B2 => n4887, C1 => n1214, C2 => 
                           n4884, A => n2077, ZN => n2076);
   U1043 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_19_port, B1 => 
                           n4878, B2 => registers_18_19_port, ZN => n2077);
   U1044 : OAI221_X1 port map( B1 => n1180, B2 => n4887, C1 => n1181, C2 => 
                           n4884, A => n2060, ZN => n2059);
   U1045 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_18_port, B1 => 
                           n4878, B2 => registers_18_18_port, ZN => n2060);
   U1046 : OAI221_X1 port map( B1 => n1147, B2 => n4887, C1 => n1148, C2 => 
                           n4884, A => n2043, ZN => n2042);
   U1047 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_17_port, B1 => 
                           n4878, B2 => registers_18_17_port, ZN => n2043);
   U1048 : OAI221_X1 port map( B1 => n1114, B2 => n4887, C1 => n1115, C2 => 
                           n4884, A => n2026, ZN => n2025);
   U1049 : AOI22_X1 port map( A1 => n4881, A2 => registers_13_16_port, B1 => 
                           n4878, B2 => registers_18_16_port, ZN => n2026);
   U1050 : OAI221_X1 port map( B1 => n4979, B2 => n1609, C1 => n4976, C2 => 
                           n1610, A => n1611, ZN => n1608);
   U1051 : AOI22_X1 port map( A1 => registers_13_31_port, A2 => n4973, B1 => 
                           registers_18_31_port, B2 => n4970, ZN => n1611);
   U1052 : OAI221_X1 port map( B1 => n4979, B2 => n1576, C1 => n4976, C2 => 
                           n1577, A => n1578, ZN => n1575);
   U1053 : AOI22_X1 port map( A1 => registers_13_30_port, A2 => n4973, B1 => 
                           registers_18_30_port, B2 => n4970, ZN => n1578);
   U1054 : OAI221_X1 port map( B1 => n4979, B2 => n1543, C1 => n4976, C2 => 
                           n1544, A => n1545, ZN => n1542);
   U1055 : AOI22_X1 port map( A1 => registers_13_29_port, A2 => n4973, B1 => 
                           registers_18_29_port, B2 => n4970, ZN => n1545);
   U1056 : OAI221_X1 port map( B1 => n4979, B2 => n1510, C1 => n4976, C2 => 
                           n1511, A => n1512, ZN => n1509);
   U1057 : AOI22_X1 port map( A1 => registers_13_28_port, A2 => n4973, B1 => 
                           registers_18_28_port, B2 => n4970, ZN => n1512);
   U1058 : OAI221_X1 port map( B1 => n4979, B2 => n1477, C1 => n4976, C2 => 
                           n1478, A => n1479, ZN => n1476);
   U1059 : AOI22_X1 port map( A1 => registers_13_27_port, A2 => n4973, B1 => 
                           registers_18_27_port, B2 => n4970, ZN => n1479);
   U1060 : OAI221_X1 port map( B1 => n4979, B2 => n1444, C1 => n4976, C2 => 
                           n1445, A => n1446, ZN => n1443);
   U1061 : AOI22_X1 port map( A1 => registers_13_26_port, A2 => n4973, B1 => 
                           registers_18_26_port, B2 => n4970, ZN => n1446);
   U1062 : OAI221_X1 port map( B1 => n4979, B2 => n1411, C1 => n4976, C2 => 
                           n1412, A => n1413, ZN => n1410);
   U1063 : AOI22_X1 port map( A1 => registers_13_25_port, A2 => n4973, B1 => 
                           registers_18_25_port, B2 => n4970, ZN => n1413);
   U1064 : OAI221_X1 port map( B1 => n4979, B2 => n1378, C1 => n4976, C2 => 
                           n1379, A => n1380, ZN => n1377);
   U1065 : AOI22_X1 port map( A1 => registers_13_24_port, A2 => n4973, B1 => 
                           registers_18_24_port, B2 => n4970, ZN => n1380);
   U1066 : OAI221_X1 port map( B1 => n4979, B2 => n1345, C1 => n4976, C2 => 
                           n1346, A => n1347, ZN => n1344);
   U1067 : AOI22_X1 port map( A1 => registers_13_23_port, A2 => n4973, B1 => 
                           registers_18_23_port, B2 => n4970, ZN => n1347);
   U1068 : OAI221_X1 port map( B1 => n4979, B2 => n1312, C1 => n4976, C2 => 
                           n1313, A => n1314, ZN => n1311);
   U1069 : AOI22_X1 port map( A1 => registers_13_22_port, A2 => n4973, B1 => 
                           registers_18_22_port, B2 => n4970, ZN => n1314);
   U1070 : OAI221_X1 port map( B1 => n4979, B2 => n1279, C1 => n4976, C2 => 
                           n1280, A => n1281, ZN => n1278);
   U1071 : AOI22_X1 port map( A1 => registers_13_21_port, A2 => n4973, B1 => 
                           registers_18_21_port, B2 => n4970, ZN => n1281);
   U1072 : OAI221_X1 port map( B1 => n4979, B2 => n1246, C1 => n4976, C2 => 
                           n1247, A => n1248, ZN => n1245);
   U1073 : AOI22_X1 port map( A1 => registers_13_20_port, A2 => n4973, B1 => 
                           registers_18_20_port, B2 => n4970, ZN => n1248);
   U1074 : OAI221_X1 port map( B1 => n4980, B2 => n1213, C1 => n4977, C2 => 
                           n1214, A => n1215, ZN => n1212);
   U1075 : AOI22_X1 port map( A1 => registers_13_19_port, A2 => n4974, B1 => 
                           registers_18_19_port, B2 => n4971, ZN => n1215);
   U1076 : OAI221_X1 port map( B1 => n4980, B2 => n1180, C1 => n4977, C2 => 
                           n1181, A => n1182, ZN => n1179);
   U1077 : AOI22_X1 port map( A1 => registers_13_18_port, A2 => n4974, B1 => 
                           registers_18_18_port, B2 => n4971, ZN => n1182);
   U1078 : OAI221_X1 port map( B1 => n4980, B2 => n1147, C1 => n4977, C2 => 
                           n1148, A => n1149, ZN => n1146);
   U1079 : AOI22_X1 port map( A1 => registers_13_17_port, A2 => n4974, B1 => 
                           registers_18_17_port, B2 => n4971, ZN => n1149);
   U1080 : OAI221_X1 port map( B1 => n4980, B2 => n1114, C1 => n4977, C2 => 
                           n1115, A => n1116, ZN => n1113);
   U1081 : AOI22_X1 port map( A1 => registers_13_16_port, A2 => n4974, B1 => 
                           registers_18_16_port, B2 => n4971, ZN => n1116);
   U1082 : OAI221_X1 port map( B1 => n4924, B2 => n833, C1 => n4921, C2 => n834
                           , A => n835, ZN => n829);
   U1083 : AOI22_X1 port map( A1 => registers_14_7_port, A2 => n4918, B1 => 
                           registers_28_7_port, B2 => n4915, ZN => n835);
   U1084 : OAI221_X1 port map( B1 => n4924, B2 => n800, C1 => n4921, C2 => n801
                           , A => n802, ZN => n796);
   U1085 : AOI22_X1 port map( A1 => registers_14_6_port, A2 => n4918, B1 => 
                           registers_28_6_port, B2 => n4915, ZN => n802);
   U1086 : OAI221_X1 port map( B1 => n4924, B2 => n767, C1 => n4921, C2 => n768
                           , A => n769, ZN => n763);
   U1087 : AOI22_X1 port map( A1 => registers_14_5_port, A2 => n4918, B1 => 
                           registers_28_5_port, B2 => n4915, ZN => n769);
   U1088 : OAI221_X1 port map( B1 => n4924, B2 => n734, C1 => n4921, C2 => n735
                           , A => n736, ZN => n730);
   U1089 : AOI22_X1 port map( A1 => registers_14_4_port, A2 => n4918, B1 => 
                           registers_28_4_port, B2 => n4915, ZN => n736);
   U1090 : OAI221_X1 port map( B1 => n4924, B2 => n701, C1 => n4921, C2 => n702
                           , A => n703, ZN => n697);
   U1091 : AOI22_X1 port map( A1 => registers_14_3_port, A2 => n4918, B1 => 
                           registers_28_3_port, B2 => n4915, ZN => n703);
   U1092 : OAI221_X1 port map( B1 => n4924, B2 => n668, C1 => n4921, C2 => n669
                           , A => n670, ZN => n664);
   U1093 : AOI22_X1 port map( A1 => registers_14_2_port, A2 => n4918, B1 => 
                           registers_28_2_port, B2 => n4915, ZN => n670);
   U1094 : OAI221_X1 port map( B1 => n4924, B2 => n635, C1 => n4921, C2 => n636
                           , A => n637, ZN => n631);
   U1095 : AOI22_X1 port map( A1 => registers_14_1_port, A2 => n4918, B1 => 
                           registers_28_1_port, B2 => n4915, ZN => n637);
   U1096 : OAI221_X1 port map( B1 => n4924, B2 => n591, C1 => n4921, C2 => n593
                           , A => n594, ZN => n584);
   U1097 : AOI22_X1 port map( A1 => registers_14_0_port, A2 => n4918, B1 => 
                           registers_28_0_port, B2 => n4915, ZN => n594);
   U1098 : OAI221_X1 port map( B1 => n833, B2 => n4831, C1 => n834, C2 => n4828
                           , A => n1879, ZN => n1877);
   U1099 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_7_port, B1 => 
                           n4820, B2 => registers_28_7_port, ZN => n1879);
   U1100 : OAI221_X1 port map( B1 => n800, B2 => n4831, C1 => n801, C2 => n4828
                           , A => n1862, ZN => n1860);
   U1101 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_6_port, B1 => 
                           n4820, B2 => registers_28_6_port, ZN => n1862);
   U1102 : OAI221_X1 port map( B1 => n767, B2 => n4831, C1 => n768, C2 => n4828
                           , A => n1845, ZN => n1834);
   U1103 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_5_port, B1 => 
                           n4820, B2 => registers_28_5_port, ZN => n1845);
   U1104 : OAI221_X1 port map( B1 => n734, B2 => n4831, C1 => n735, C2 => n4828
                           , A => n1764, ZN => n1762);
   U1105 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_4_port, B1 => 
                           n4820, B2 => registers_28_4_port, ZN => n1764);
   U1106 : OAI221_X1 port map( B1 => n701, B2 => n4831, C1 => n702, C2 => n4828
                           , A => n1747, ZN => n1745);
   U1107 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_3_port, B1 => 
                           n4820, B2 => registers_28_3_port, ZN => n1747);
   U1108 : OAI221_X1 port map( B1 => n668, B2 => n4831, C1 => n669, C2 => n4828
                           , A => n1730, ZN => n1728);
   U1109 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_2_port, B1 => 
                           n4820, B2 => registers_28_2_port, ZN => n1730);
   U1110 : OAI221_X1 port map( B1 => n635, B2 => n4831, C1 => n636, C2 => n4828
                           , A => n1713, ZN => n1711);
   U1111 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_1_port, B1 => 
                           n4820, B2 => registers_28_1_port, ZN => n1713);
   U1112 : OAI221_X1 port map( B1 => n591, B2 => n4831, C1 => n593, C2 => n4828
                           , A => n1686, ZN => n1680);
   U1113 : AOI22_X1 port map( A1 => n4825, A2 => registers_14_0_port, B1 => 
                           n4820, B2 => registers_28_0_port, ZN => n1686);
   U1114 : OAI221_X1 port map( B1 => n1097, B2 => n4830, C1 => n1098, C2 => 
                           n4827, A => n2015, ZN => n2013);
   U1115 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_15_port, B1 => 
                           n4821, B2 => registers_28_15_port, ZN => n2015);
   U1116 : OAI221_X1 port map( B1 => n1064, B2 => n4830, C1 => n1065, C2 => 
                           n4827, A => n1998, ZN => n1996);
   U1117 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_14_port, B1 => 
                           n4821, B2 => registers_28_14_port, ZN => n1998);
   U1118 : OAI221_X1 port map( B1 => n1031, B2 => n4830, C1 => n1032, C2 => 
                           n4827, A => n1981, ZN => n1979);
   U1119 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_13_port, B1 => 
                           n4821, B2 => registers_28_13_port, ZN => n1981);
   U1120 : OAI221_X1 port map( B1 => n998, B2 => n4830, C1 => n999, C2 => n4827
                           , A => n1964, ZN => n1962);
   U1121 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_12_port, B1 => 
                           n4821, B2 => registers_28_12_port, ZN => n1964);
   U1122 : OAI221_X1 port map( B1 => n965, B2 => n4830, C1 => n966, C2 => n4827
                           , A => n1947, ZN => n1945);
   U1123 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_11_port, B1 => 
                           n4820, B2 => registers_28_11_port, ZN => n1947);
   U1124 : OAI221_X1 port map( B1 => n932, B2 => n4830, C1 => n933, C2 => n4827
                           , A => n1930, ZN => n1928);
   U1125 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_10_port, B1 => 
                           n4820, B2 => registers_28_10_port, ZN => n1930);
   U1126 : OAI221_X1 port map( B1 => n899, B2 => n4830, C1 => n900, C2 => n4827
                           , A => n1913, ZN => n1911);
   U1127 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_9_port, B1 => 
                           n4820, B2 => registers_28_9_port, ZN => n1913);
   U1128 : OAI221_X1 port map( B1 => n866, B2 => n4830, C1 => n867, C2 => n4827
                           , A => n1896, ZN => n1894);
   U1129 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_8_port, B1 => 
                           n4820, B2 => registers_28_8_port, ZN => n1896);
   U1130 : OAI221_X1 port map( B1 => n4923, B2 => n1097, C1 => n4920, C2 => 
                           n1098, A => n1099, ZN => n1093);
   U1131 : AOI22_X1 port map( A1 => registers_14_15_port, A2 => n4917, B1 => 
                           registers_28_15_port, B2 => n4914, ZN => n1099);
   U1132 : OAI221_X1 port map( B1 => n4923, B2 => n1064, C1 => n4920, C2 => 
                           n1065, A => n1066, ZN => n1060);
   U1133 : AOI22_X1 port map( A1 => registers_14_14_port, A2 => n4917, B1 => 
                           registers_28_14_port, B2 => n4914, ZN => n1066);
   U1134 : OAI221_X1 port map( B1 => n4923, B2 => n1031, C1 => n4920, C2 => 
                           n1032, A => n1033, ZN => n1027);
   U1135 : AOI22_X1 port map( A1 => registers_14_13_port, A2 => n4917, B1 => 
                           registers_28_13_port, B2 => n4914, ZN => n1033);
   U1136 : OAI221_X1 port map( B1 => n4923, B2 => n998, C1 => n4920, C2 => n999
                           , A => n1000, ZN => n994);
   U1137 : AOI22_X1 port map( A1 => registers_14_12_port, A2 => n4917, B1 => 
                           registers_28_12_port, B2 => n4914, ZN => n1000);
   U1138 : OAI221_X1 port map( B1 => n4923, B2 => n965, C1 => n4920, C2 => n966
                           , A => n967, ZN => n961);
   U1139 : AOI22_X1 port map( A1 => registers_14_11_port, A2 => n4917, B1 => 
                           registers_28_11_port, B2 => n4914, ZN => n967);
   U1140 : OAI221_X1 port map( B1 => n4923, B2 => n932, C1 => n4920, C2 => n933
                           , A => n934, ZN => n928);
   U1141 : AOI22_X1 port map( A1 => registers_14_10_port, A2 => n4917, B1 => 
                           registers_28_10_port, B2 => n4914, ZN => n934);
   U1142 : OAI221_X1 port map( B1 => n4923, B2 => n899, C1 => n4920, C2 => n900
                           , A => n901, ZN => n895);
   U1143 : AOI22_X1 port map( A1 => registers_14_9_port, A2 => n4917, B1 => 
                           registers_28_9_port, B2 => n4914, ZN => n901);
   U1144 : OAI221_X1 port map( B1 => n4923, B2 => n866, C1 => n4920, C2 => n867
                           , A => n868, ZN => n862);
   U1145 : AOI22_X1 port map( A1 => registers_14_8_port, A2 => n4917, B1 => 
                           registers_28_8_port, B2 => n4914, ZN => n868);
   U1146 : OAI221_X1 port map( B1 => n1638, B2 => n4829, C1 => n1639, C2 => 
                           n4826, A => n2300, ZN => n2297);
   U1147 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_31_port, B1 => 
                           n4822, B2 => registers_28_31_port, ZN => n2300);
   U1148 : OAI221_X1 port map( B1 => n1592, B2 => n4829, C1 => n1593, C2 => 
                           n4826, A => n2270, ZN => n2268);
   U1149 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_30_port, B1 => 
                           n4822, B2 => registers_28_30_port, ZN => n2270);
   U1150 : OAI221_X1 port map( B1 => n1559, B2 => n4829, C1 => n1560, C2 => 
                           n4826, A => n2253, ZN => n2251);
   U1151 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_29_port, B1 => 
                           n4822, B2 => registers_28_29_port, ZN => n2253);
   U1152 : OAI221_X1 port map( B1 => n1526, B2 => n4829, C1 => n1527, C2 => 
                           n4826, A => n2236, ZN => n2234);
   U1153 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_28_port, B1 => 
                           n4822, B2 => registers_28_28_port, ZN => n2236);
   U1154 : OAI221_X1 port map( B1 => n1493, B2 => n4829, C1 => n1494, C2 => 
                           n4826, A => n2219, ZN => n2217);
   U1155 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_27_port, B1 => 
                           n4822, B2 => registers_28_27_port, ZN => n2219);
   U1156 : OAI221_X1 port map( B1 => n1460, B2 => n4829, C1 => n1461, C2 => 
                           n4826, A => n2202, ZN => n2200);
   U1157 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_26_port, B1 => 
                           n4822, B2 => registers_28_26_port, ZN => n2202);
   U1158 : OAI221_X1 port map( B1 => n1427, B2 => n4829, C1 => n1428, C2 => 
                           n4826, A => n2185, ZN => n2183);
   U1159 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_25_port, B1 => 
                           n4822, B2 => registers_28_25_port, ZN => n2185);
   U1160 : OAI221_X1 port map( B1 => n1394, B2 => n4829, C1 => n1395, C2 => 
                           n4826, A => n2168, ZN => n2166);
   U1161 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_24_port, B1 => 
                           n4822, B2 => registers_28_24_port, ZN => n2168);
   U1162 : OAI221_X1 port map( B1 => n1361, B2 => n4829, C1 => n1362, C2 => 
                           n4826, A => n2151, ZN => n2149);
   U1163 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_23_port, B1 => 
                           n4821, B2 => registers_28_23_port, ZN => n2151);
   U1164 : OAI221_X1 port map( B1 => n1328, B2 => n4829, C1 => n1329, C2 => 
                           n4826, A => n2134, ZN => n2132);
   U1165 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_22_port, B1 => 
                           n4821, B2 => registers_28_22_port, ZN => n2134);
   U1166 : OAI221_X1 port map( B1 => n1295, B2 => n4829, C1 => n1296, C2 => 
                           n4826, A => n2117, ZN => n2115);
   U1167 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_21_port, B1 => 
                           n4821, B2 => registers_28_21_port, ZN => n2117);
   U1168 : OAI221_X1 port map( B1 => n1262, B2 => n4829, C1 => n1263, C2 => 
                           n4826, A => n2100, ZN => n2098);
   U1169 : AOI22_X1 port map( A1 => n4823, A2 => registers_14_20_port, B1 => 
                           n4821, B2 => registers_28_20_port, ZN => n2100);
   U1170 : OAI221_X1 port map( B1 => n1229, B2 => n4830, C1 => n1230, C2 => 
                           n4827, A => n2083, ZN => n2081);
   U1171 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_19_port, B1 => 
                           n4821, B2 => registers_28_19_port, ZN => n2083);
   U1172 : OAI221_X1 port map( B1 => n1196, B2 => n4830, C1 => n1197, C2 => 
                           n4827, A => n2066, ZN => n2064);
   U1173 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_18_port, B1 => 
                           n4821, B2 => registers_28_18_port, ZN => n2066);
   U1174 : OAI221_X1 port map( B1 => n1163, B2 => n4830, C1 => n1164, C2 => 
                           n4827, A => n2049, ZN => n2047);
   U1175 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_17_port, B1 => 
                           n4821, B2 => registers_28_17_port, ZN => n2049);
   U1176 : OAI221_X1 port map( B1 => n1130, B2 => n4830, C1 => n1131, C2 => 
                           n4827, A => n2032, ZN => n2030);
   U1177 : AOI22_X1 port map( A1 => n4824, A2 => registers_14_16_port, B1 => 
                           n4821, B2 => registers_28_16_port, ZN => n2032);
   U1178 : OAI221_X1 port map( B1 => n4922, B2 => n1638, C1 => n4919, C2 => 
                           n1639, A => n1640, ZN => n1633);
   U1179 : AOI22_X1 port map( A1 => registers_14_31_port, A2 => n4916, B1 => 
                           registers_28_31_port, B2 => n4913, ZN => n1640);
   U1180 : OAI221_X1 port map( B1 => n4922, B2 => n1592, C1 => n4919, C2 => 
                           n1593, A => n1594, ZN => n1588);
   U1181 : AOI22_X1 port map( A1 => registers_14_30_port, A2 => n4916, B1 => 
                           registers_28_30_port, B2 => n4913, ZN => n1594);
   U1182 : OAI221_X1 port map( B1 => n4922, B2 => n1559, C1 => n4919, C2 => 
                           n1560, A => n1561, ZN => n1555);
   U1183 : AOI22_X1 port map( A1 => registers_14_29_port, A2 => n4916, B1 => 
                           registers_28_29_port, B2 => n4913, ZN => n1561);
   U1184 : OAI221_X1 port map( B1 => n4922, B2 => n1526, C1 => n4919, C2 => 
                           n1527, A => n1528, ZN => n1522);
   U1185 : AOI22_X1 port map( A1 => registers_14_28_port, A2 => n4916, B1 => 
                           registers_28_28_port, B2 => n4913, ZN => n1528);
   U1186 : OAI221_X1 port map( B1 => n4922, B2 => n1493, C1 => n4919, C2 => 
                           n1494, A => n1495, ZN => n1489);
   U1187 : AOI22_X1 port map( A1 => registers_14_27_port, A2 => n4916, B1 => 
                           registers_28_27_port, B2 => n4913, ZN => n1495);
   U1188 : OAI221_X1 port map( B1 => n4922, B2 => n1460, C1 => n4919, C2 => 
                           n1461, A => n1462, ZN => n1456);
   U1189 : AOI22_X1 port map( A1 => registers_14_26_port, A2 => n4916, B1 => 
                           registers_28_26_port, B2 => n4913, ZN => n1462);
   U1190 : OAI221_X1 port map( B1 => n4922, B2 => n1427, C1 => n4919, C2 => 
                           n1428, A => n1429, ZN => n1423);
   U1191 : AOI22_X1 port map( A1 => registers_14_25_port, A2 => n4916, B1 => 
                           registers_28_25_port, B2 => n4913, ZN => n1429);
   U1192 : OAI221_X1 port map( B1 => n4922, B2 => n1394, C1 => n4919, C2 => 
                           n1395, A => n1396, ZN => n1390);
   U1193 : AOI22_X1 port map( A1 => registers_14_24_port, A2 => n4916, B1 => 
                           registers_28_24_port, B2 => n4913, ZN => n1396);
   U1194 : OAI221_X1 port map( B1 => n4922, B2 => n1361, C1 => n4919, C2 => 
                           n1362, A => n1363, ZN => n1357);
   U1195 : AOI22_X1 port map( A1 => registers_14_23_port, A2 => n4916, B1 => 
                           registers_28_23_port, B2 => n4913, ZN => n1363);
   U1196 : OAI221_X1 port map( B1 => n4922, B2 => n1328, C1 => n4919, C2 => 
                           n1329, A => n1330, ZN => n1324);
   U1197 : AOI22_X1 port map( A1 => registers_14_22_port, A2 => n4916, B1 => 
                           registers_28_22_port, B2 => n4913, ZN => n1330);
   U1198 : OAI221_X1 port map( B1 => n4922, B2 => n1295, C1 => n4919, C2 => 
                           n1296, A => n1297, ZN => n1291);
   U1199 : AOI22_X1 port map( A1 => registers_14_21_port, A2 => n4916, B1 => 
                           registers_28_21_port, B2 => n4913, ZN => n1297);
   U1200 : OAI221_X1 port map( B1 => n4922, B2 => n1262, C1 => n4919, C2 => 
                           n1263, A => n1264, ZN => n1258);
   U1201 : AOI22_X1 port map( A1 => registers_14_20_port, A2 => n4916, B1 => 
                           registers_28_20_port, B2 => n4913, ZN => n1264);
   U1202 : OAI221_X1 port map( B1 => n4923, B2 => n1229, C1 => n4920, C2 => 
                           n1230, A => n1231, ZN => n1225);
   U1203 : AOI22_X1 port map( A1 => registers_14_19_port, A2 => n4917, B1 => 
                           registers_28_19_port, B2 => n4914, ZN => n1231);
   U1204 : OAI221_X1 port map( B1 => n4923, B2 => n1196, C1 => n4920, C2 => 
                           n1197, A => n1198, ZN => n1192);
   U1205 : AOI22_X1 port map( A1 => registers_14_18_port, A2 => n4917, B1 => 
                           registers_28_18_port, B2 => n4914, ZN => n1198);
   U1206 : OAI221_X1 port map( B1 => n4923, B2 => n1163, C1 => n4920, C2 => 
                           n1164, A => n1165, ZN => n1159);
   U1207 : AOI22_X1 port map( A1 => registers_14_17_port, A2 => n4917, B1 => 
                           registers_28_17_port, B2 => n4914, ZN => n1165);
   U1208 : OAI221_X1 port map( B1 => n4923, B2 => n1130, C1 => n4920, C2 => 
                           n1131, A => n1132, ZN => n1126);
   U1209 : AOI22_X1 port map( A1 => registers_14_16_port, A2 => n4917, B1 => 
                           registers_28_16_port, B2 => n4914, ZN => n1132);
   U1210 : AOI22_X1 port map( A1 => registers_12_7_port, A2 => n4963, B1 => 
                           registers_30_7_port, B2 => n4960, ZN => n822);
   U1211 : AOI22_X1 port map( A1 => registers_20_7_port, A2 => n4951, B1 => 
                           registers_21_7_port, B2 => n4948, ZN => n825);
   U1212 : AOI22_X1 port map( A1 => registers_24_7_port, A2 => n4939, B1 => 
                           registers_25_7_port, B2 => n4936, ZN => n828);
   U1213 : AOI22_X1 port map( A1 => registers_12_6_port, A2 => n4963, B1 => 
                           registers_30_6_port, B2 => n4960, ZN => n789);
   U1214 : AOI22_X1 port map( A1 => registers_20_6_port, A2 => n4951, B1 => 
                           registers_21_6_port, B2 => n4948, ZN => n792);
   U1215 : AOI22_X1 port map( A1 => registers_24_6_port, A2 => n4939, B1 => 
                           registers_25_6_port, B2 => n4936, ZN => n795);
   U1216 : AOI22_X1 port map( A1 => registers_12_5_port, A2 => n4963, B1 => 
                           registers_30_5_port, B2 => n4960, ZN => n756);
   U1217 : AOI22_X1 port map( A1 => registers_20_5_port, A2 => n4951, B1 => 
                           registers_21_5_port, B2 => n4948, ZN => n759);
   U1218 : AOI22_X1 port map( A1 => registers_24_5_port, A2 => n4939, B1 => 
                           registers_25_5_port, B2 => n4936, ZN => n762);
   U1219 : AOI22_X1 port map( A1 => registers_12_4_port, A2 => n4963, B1 => 
                           registers_30_4_port, B2 => n4960, ZN => n723);
   U1220 : AOI22_X1 port map( A1 => registers_20_4_port, A2 => n4951, B1 => 
                           registers_21_4_port, B2 => n4948, ZN => n726);
   U1221 : AOI22_X1 port map( A1 => registers_24_4_port, A2 => n4939, B1 => 
                           registers_25_4_port, B2 => n4936, ZN => n729);
   U1222 : AOI22_X1 port map( A1 => registers_12_3_port, A2 => n4963, B1 => 
                           registers_30_3_port, B2 => n4960, ZN => n690);
   U1223 : AOI22_X1 port map( A1 => registers_20_3_port, A2 => n4951, B1 => 
                           registers_21_3_port, B2 => n4948, ZN => n693);
   U1224 : AOI22_X1 port map( A1 => registers_24_3_port, A2 => n4939, B1 => 
                           registers_25_3_port, B2 => n4936, ZN => n696);
   U1225 : AOI22_X1 port map( A1 => registers_12_2_port, A2 => n4963, B1 => 
                           registers_30_2_port, B2 => n4960, ZN => n657);
   U1226 : AOI22_X1 port map( A1 => registers_20_2_port, A2 => n4951, B1 => 
                           registers_21_2_port, B2 => n4948, ZN => n660);
   U1227 : AOI22_X1 port map( A1 => registers_24_2_port, A2 => n4939, B1 => 
                           registers_25_2_port, B2 => n4936, ZN => n663);
   U1228 : AOI22_X1 port map( A1 => registers_12_1_port, A2 => n4963, B1 => 
                           registers_30_1_port, B2 => n4960, ZN => n624);
   U1229 : AOI22_X1 port map( A1 => registers_20_1_port, A2 => n4951, B1 => 
                           registers_21_1_port, B2 => n4948, ZN => n627);
   U1230 : AOI22_X1 port map( A1 => registers_24_1_port, A2 => n4939, B1 => 
                           registers_25_1_port, B2 => n4936, ZN => n630);
   U1231 : AOI22_X1 port map( A1 => registers_12_0_port, A2 => n4963, B1 => 
                           registers_30_0_port, B2 => n4960, ZN => n566);
   U1232 : AOI22_X1 port map( A1 => registers_20_0_port, A2 => n4951, B1 => 
                           registers_21_0_port, B2 => n4948, ZN => n573);
   U1233 : AOI22_X1 port map( A1 => registers_24_0_port, A2 => n4939, B1 => 
                           registers_25_0_port, B2 => n4936, ZN => n580);
   U1234 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_15_port, B1 => 
                           n4866, B2 => registers_30_15_port, ZN => n2010);
   U1235 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_15_port, B1 => 
                           n4854, B2 => registers_21_15_port, ZN => n2011);
   U1236 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_15_port, B1 => 
                           n4842, B2 => registers_25_15_port, ZN => n2012);
   U1237 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_14_port, B1 => 
                           n4866, B2 => registers_30_14_port, ZN => n1993);
   U1238 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_14_port, B1 => 
                           n4854, B2 => registers_21_14_port, ZN => n1994);
   U1239 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_14_port, B1 => 
                           n4842, B2 => registers_25_14_port, ZN => n1995);
   U1240 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_13_port, B1 => 
                           n4866, B2 => registers_30_13_port, ZN => n1976);
   U1241 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_13_port, B1 => 
                           n4854, B2 => registers_21_13_port, ZN => n1977);
   U1242 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_13_port, B1 => 
                           n4842, B2 => registers_25_13_port, ZN => n1978);
   U1243 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_12_port, B1 => 
                           n4866, B2 => registers_30_12_port, ZN => n1959);
   U1244 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_12_port, B1 => 
                           n4854, B2 => registers_21_12_port, ZN => n1960);
   U1245 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_12_port, B1 => 
                           n4842, B2 => registers_25_12_port, ZN => n1961);
   U1246 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_11_port, B1 => 
                           n4865, B2 => registers_30_11_port, ZN => n1942);
   U1247 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_11_port, B1 => 
                           n4853, B2 => registers_21_11_port, ZN => n1943);
   U1248 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_11_port, B1 => 
                           n4841, B2 => registers_25_11_port, ZN => n1944);
   U1249 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_10_port, B1 => 
                           n4865, B2 => registers_30_10_port, ZN => n1925);
   U1250 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_10_port, B1 => 
                           n4853, B2 => registers_21_10_port, ZN => n1926);
   U1251 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_10_port, B1 => 
                           n4841, B2 => registers_25_10_port, ZN => n1927);
   U1252 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_9_port, B1 => 
                           n4865, B2 => registers_30_9_port, ZN => n1908);
   U1253 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_9_port, B1 => 
                           n4853, B2 => registers_21_9_port, ZN => n1909);
   U1254 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_9_port, B1 => 
                           n4841, B2 => registers_25_9_port, ZN => n1910);
   U1255 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_8_port, B1 => 
                           n4865, B2 => registers_30_8_port, ZN => n1891);
   U1256 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_8_port, B1 => 
                           n4853, B2 => registers_21_8_port, ZN => n1892);
   U1257 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_8_port, B1 => 
                           n4841, B2 => registers_25_8_port, ZN => n1893);
   U1258 : AOI22_X1 port map( A1 => registers_12_15_port, A2 => n4962, B1 => 
                           registers_30_15_port, B2 => n4959, ZN => n1086);
   U1259 : AOI22_X1 port map( A1 => registers_20_15_port, A2 => n4950, B1 => 
                           registers_21_15_port, B2 => n4947, ZN => n1089);
   U1260 : AOI22_X1 port map( A1 => registers_24_15_port, A2 => n4938, B1 => 
                           registers_25_15_port, B2 => n4935, ZN => n1092);
   U1261 : AOI22_X1 port map( A1 => registers_12_14_port, A2 => n4962, B1 => 
                           registers_30_14_port, B2 => n4959, ZN => n1053);
   U1262 : AOI22_X1 port map( A1 => registers_20_14_port, A2 => n4950, B1 => 
                           registers_21_14_port, B2 => n4947, ZN => n1056);
   U1263 : AOI22_X1 port map( A1 => registers_24_14_port, A2 => n4938, B1 => 
                           registers_25_14_port, B2 => n4935, ZN => n1059);
   U1264 : AOI22_X1 port map( A1 => registers_12_13_port, A2 => n4962, B1 => 
                           registers_30_13_port, B2 => n4959, ZN => n1020);
   U1265 : AOI22_X1 port map( A1 => registers_20_13_port, A2 => n4950, B1 => 
                           registers_21_13_port, B2 => n4947, ZN => n1023);
   U1266 : AOI22_X1 port map( A1 => registers_24_13_port, A2 => n4938, B1 => 
                           registers_25_13_port, B2 => n4935, ZN => n1026);
   U1267 : AOI22_X1 port map( A1 => registers_12_12_port, A2 => n4962, B1 => 
                           registers_30_12_port, B2 => n4959, ZN => n987);
   U1268 : AOI22_X1 port map( A1 => registers_20_12_port, A2 => n4950, B1 => 
                           registers_21_12_port, B2 => n4947, ZN => n990);
   U1269 : AOI22_X1 port map( A1 => registers_24_12_port, A2 => n4938, B1 => 
                           registers_25_12_port, B2 => n4935, ZN => n993);
   U1270 : AOI22_X1 port map( A1 => registers_12_11_port, A2 => n4962, B1 => 
                           registers_30_11_port, B2 => n4959, ZN => n954);
   U1271 : AOI22_X1 port map( A1 => registers_20_11_port, A2 => n4950, B1 => 
                           registers_21_11_port, B2 => n4947, ZN => n957);
   U1272 : AOI22_X1 port map( A1 => registers_24_11_port, A2 => n4938, B1 => 
                           registers_25_11_port, B2 => n4935, ZN => n960);
   U1273 : AOI22_X1 port map( A1 => registers_12_10_port, A2 => n4962, B1 => 
                           registers_30_10_port, B2 => n4959, ZN => n921);
   U1274 : AOI22_X1 port map( A1 => registers_20_10_port, A2 => n4950, B1 => 
                           registers_21_10_port, B2 => n4947, ZN => n924);
   U1275 : AOI22_X1 port map( A1 => registers_24_10_port, A2 => n4938, B1 => 
                           registers_25_10_port, B2 => n4935, ZN => n927);
   U1276 : AOI22_X1 port map( A1 => registers_12_9_port, A2 => n4962, B1 => 
                           registers_30_9_port, B2 => n4959, ZN => n888);
   U1277 : AOI22_X1 port map( A1 => registers_20_9_port, A2 => n4950, B1 => 
                           registers_21_9_port, B2 => n4947, ZN => n891);
   U1278 : AOI22_X1 port map( A1 => registers_24_9_port, A2 => n4938, B1 => 
                           registers_25_9_port, B2 => n4935, ZN => n894);
   U1279 : AOI22_X1 port map( A1 => registers_12_8_port, A2 => n4962, B1 => 
                           registers_30_8_port, B2 => n4959, ZN => n855);
   U1280 : AOI22_X1 port map( A1 => registers_20_8_port, A2 => n4950, B1 => 
                           registers_21_8_port, B2 => n4947, ZN => n858);
   U1281 : AOI22_X1 port map( A1 => registers_24_8_port, A2 => n4938, B1 => 
                           registers_25_8_port, B2 => n4935, ZN => n861);
   U1282 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_7_port, B1 => 
                           n4865, B2 => registers_30_7_port, ZN => n1874);
   U1283 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_7_port, B1 => 
                           n4853, B2 => registers_21_7_port, ZN => n1875);
   U1284 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_7_port, B1 => 
                           n4841, B2 => registers_25_7_port, ZN => n1876);
   U1285 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_6_port, B1 => 
                           n4865, B2 => registers_30_6_port, ZN => n1857);
   U1286 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_6_port, B1 => 
                           n4853, B2 => registers_21_6_port, ZN => n1858);
   U1287 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_6_port, B1 => 
                           n4841, B2 => registers_25_6_port, ZN => n1859);
   U1288 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_5_port, B1 => 
                           n4865, B2 => registers_30_5_port, ZN => n1776);
   U1289 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_5_port, B1 => 
                           n4853, B2 => registers_21_5_port, ZN => n1777);
   U1290 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_5_port, B1 => 
                           n4841, B2 => registers_25_5_port, ZN => n1801);
   U1291 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_4_port, B1 => 
                           n4865, B2 => registers_30_4_port, ZN => n1759);
   U1292 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_4_port, B1 => 
                           n4853, B2 => registers_21_4_port, ZN => n1760);
   U1293 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_4_port, B1 => 
                           n4841, B2 => registers_25_4_port, ZN => n1761);
   U1294 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_3_port, B1 => 
                           n4865, B2 => registers_30_3_port, ZN => n1742);
   U1295 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_3_port, B1 => 
                           n4853, B2 => registers_21_3_port, ZN => n1743);
   U1296 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_3_port, B1 => 
                           n4841, B2 => registers_25_3_port, ZN => n1744);
   U1297 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_2_port, B1 => 
                           n4865, B2 => registers_30_2_port, ZN => n1725);
   U1298 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_2_port, B1 => 
                           n4853, B2 => registers_21_2_port, ZN => n1726);
   U1299 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_2_port, B1 => 
                           n4841, B2 => registers_25_2_port, ZN => n1727);
   U1300 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_1_port, B1 => 
                           n4865, B2 => registers_30_1_port, ZN => n1708);
   U1301 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_1_port, B1 => 
                           n4853, B2 => registers_21_1_port, ZN => n1709);
   U1302 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_1_port, B1 => 
                           n4841, B2 => registers_25_1_port, ZN => n1710);
   U1303 : AOI22_X1 port map( A1 => n4870, A2 => registers_12_0_port, B1 => 
                           n4865, B2 => registers_30_0_port, ZN => n1666);
   U1304 : AOI22_X1 port map( A1 => n4858, A2 => registers_20_0_port, B1 => 
                           n4853, B2 => registers_21_0_port, ZN => n1671);
   U1305 : AOI22_X1 port map( A1 => n4846, A2 => registers_24_0_port, B1 => 
                           n4841, B2 => registers_25_0_port, ZN => n1676);
   U1306 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_31_port, B1 => 
                           n4867, B2 => registers_30_31_port, ZN => n2289);
   U1307 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_31_port, B1 => 
                           n4855, B2 => registers_21_31_port, ZN => n2293);
   U1308 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_31_port, B1 => 
                           n4843, B2 => registers_25_31_port, ZN => n2296);
   U1309 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_30_port, B1 => 
                           n4867, B2 => registers_30_30_port, ZN => n2265);
   U1310 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_30_port, B1 => 
                           n4855, B2 => registers_21_30_port, ZN => n2266);
   U1311 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_30_port, B1 => 
                           n4843, B2 => registers_25_30_port, ZN => n2267);
   U1312 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_29_port, B1 => 
                           n4867, B2 => registers_30_29_port, ZN => n2248);
   U1313 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_29_port, B1 => 
                           n4855, B2 => registers_21_29_port, ZN => n2249);
   U1314 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_29_port, B1 => 
                           n4843, B2 => registers_25_29_port, ZN => n2250);
   U1315 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_28_port, B1 => 
                           n4867, B2 => registers_30_28_port, ZN => n2231);
   U1316 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_28_port, B1 => 
                           n4855, B2 => registers_21_28_port, ZN => n2232);
   U1317 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_28_port, B1 => 
                           n4843, B2 => registers_25_28_port, ZN => n2233);
   U1318 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_27_port, B1 => 
                           n4867, B2 => registers_30_27_port, ZN => n2214);
   U1319 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_27_port, B1 => 
                           n4855, B2 => registers_21_27_port, ZN => n2215);
   U1320 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_27_port, B1 => 
                           n4843, B2 => registers_25_27_port, ZN => n2216);
   U1321 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_26_port, B1 => 
                           n4867, B2 => registers_30_26_port, ZN => n2197);
   U1322 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_26_port, B1 => 
                           n4855, B2 => registers_21_26_port, ZN => n2198);
   U1323 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_26_port, B1 => 
                           n4843, B2 => registers_25_26_port, ZN => n2199);
   U1324 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_25_port, B1 => 
                           n4867, B2 => registers_30_25_port, ZN => n2180);
   U1325 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_25_port, B1 => 
                           n4855, B2 => registers_21_25_port, ZN => n2181);
   U1326 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_25_port, B1 => 
                           n4843, B2 => registers_25_25_port, ZN => n2182);
   U1327 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_24_port, B1 => 
                           n4867, B2 => registers_30_24_port, ZN => n2163);
   U1328 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_24_port, B1 => 
                           n4855, B2 => registers_21_24_port, ZN => n2164);
   U1329 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_24_port, B1 => 
                           n4843, B2 => registers_25_24_port, ZN => n2165);
   U1330 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_23_port, B1 => 
                           n4866, B2 => registers_30_23_port, ZN => n2146);
   U1331 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_23_port, B1 => 
                           n4854, B2 => registers_21_23_port, ZN => n2147);
   U1332 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_23_port, B1 => 
                           n4842, B2 => registers_25_23_port, ZN => n2148);
   U1333 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_22_port, B1 => 
                           n4866, B2 => registers_30_22_port, ZN => n2129);
   U1334 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_22_port, B1 => 
                           n4854, B2 => registers_21_22_port, ZN => n2130);
   U1335 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_22_port, B1 => 
                           n4842, B2 => registers_25_22_port, ZN => n2131);
   U1336 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_21_port, B1 => 
                           n4866, B2 => registers_30_21_port, ZN => n2112);
   U1337 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_21_port, B1 => 
                           n4854, B2 => registers_21_21_port, ZN => n2113);
   U1338 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_21_port, B1 => 
                           n4842, B2 => registers_25_21_port, ZN => n2114);
   U1339 : AOI22_X1 port map( A1 => n4868, A2 => registers_12_20_port, B1 => 
                           n4866, B2 => registers_30_20_port, ZN => n2095);
   U1340 : AOI22_X1 port map( A1 => n4856, A2 => registers_20_20_port, B1 => 
                           n4854, B2 => registers_21_20_port, ZN => n2096);
   U1341 : AOI22_X1 port map( A1 => n4844, A2 => registers_24_20_port, B1 => 
                           n4842, B2 => registers_25_20_port, ZN => n2097);
   U1342 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_19_port, B1 => 
                           n4866, B2 => registers_30_19_port, ZN => n2078);
   U1343 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_19_port, B1 => 
                           n4854, B2 => registers_21_19_port, ZN => n2079);
   U1344 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_19_port, B1 => 
                           n4842, B2 => registers_25_19_port, ZN => n2080);
   U1345 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_18_port, B1 => 
                           n4866, B2 => registers_30_18_port, ZN => n2061);
   U1346 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_18_port, B1 => 
                           n4854, B2 => registers_21_18_port, ZN => n2062);
   U1347 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_18_port, B1 => 
                           n4842, B2 => registers_25_18_port, ZN => n2063);
   U1348 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_17_port, B1 => 
                           n4866, B2 => registers_30_17_port, ZN => n2044);
   U1349 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_17_port, B1 => 
                           n4854, B2 => registers_21_17_port, ZN => n2045);
   U1350 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_17_port, B1 => 
                           n4842, B2 => registers_25_17_port, ZN => n2046);
   U1351 : AOI22_X1 port map( A1 => n4869, A2 => registers_12_16_port, B1 => 
                           n4866, B2 => registers_30_16_port, ZN => n2027);
   U1352 : AOI22_X1 port map( A1 => n4857, A2 => registers_20_16_port, B1 => 
                           n4854, B2 => registers_21_16_port, ZN => n2028);
   U1353 : AOI22_X1 port map( A1 => n4845, A2 => registers_24_16_port, B1 => 
                           n4842, B2 => registers_25_16_port, ZN => n2029);
   U1354 : AOI22_X1 port map( A1 => registers_12_31_port, A2 => n4961, B1 => 
                           registers_30_31_port, B2 => n4958, ZN => n1621);
   U1355 : AOI22_X1 port map( A1 => registers_20_31_port, A2 => n4949, B1 => 
                           registers_21_31_port, B2 => n4946, ZN => n1627);
   U1356 : AOI22_X1 port map( A1 => registers_24_31_port, A2 => n4937, B1 => 
                           registers_25_31_port, B2 => n4934, ZN => n1632);
   U1357 : AOI22_X1 port map( A1 => registers_12_30_port, A2 => n4961, B1 => 
                           registers_30_30_port, B2 => n4958, ZN => n1581);
   U1358 : AOI22_X1 port map( A1 => registers_20_30_port, A2 => n4949, B1 => 
                           registers_21_30_port, B2 => n4946, ZN => n1584);
   U1359 : AOI22_X1 port map( A1 => registers_24_30_port, A2 => n4937, B1 => 
                           registers_25_30_port, B2 => n4934, ZN => n1587);
   U1360 : AOI22_X1 port map( A1 => registers_12_29_port, A2 => n4961, B1 => 
                           registers_30_29_port, B2 => n4958, ZN => n1548);
   U1361 : AOI22_X1 port map( A1 => registers_20_29_port, A2 => n4949, B1 => 
                           registers_21_29_port, B2 => n4946, ZN => n1551);
   U1362 : AOI22_X1 port map( A1 => registers_24_29_port, A2 => n4937, B1 => 
                           registers_25_29_port, B2 => n4934, ZN => n1554);
   U1363 : AOI22_X1 port map( A1 => registers_12_28_port, A2 => n4961, B1 => 
                           registers_30_28_port, B2 => n4958, ZN => n1515);
   U1364 : AOI22_X1 port map( A1 => registers_20_28_port, A2 => n4949, B1 => 
                           registers_21_28_port, B2 => n4946, ZN => n1518);
   U1365 : AOI22_X1 port map( A1 => registers_24_28_port, A2 => n4937, B1 => 
                           registers_25_28_port, B2 => n4934, ZN => n1521);
   U1366 : AOI22_X1 port map( A1 => registers_12_27_port, A2 => n4961, B1 => 
                           registers_30_27_port, B2 => n4958, ZN => n1482);
   U1367 : AOI22_X1 port map( A1 => registers_20_27_port, A2 => n4949, B1 => 
                           registers_21_27_port, B2 => n4946, ZN => n1485);
   U1368 : AOI22_X1 port map( A1 => registers_24_27_port, A2 => n4937, B1 => 
                           registers_25_27_port, B2 => n4934, ZN => n1488);
   U1369 : AOI22_X1 port map( A1 => registers_12_26_port, A2 => n4961, B1 => 
                           registers_30_26_port, B2 => n4958, ZN => n1449);
   U1370 : AOI22_X1 port map( A1 => registers_20_26_port, A2 => n4949, B1 => 
                           registers_21_26_port, B2 => n4946, ZN => n1452);
   U1371 : AOI22_X1 port map( A1 => registers_24_26_port, A2 => n4937, B1 => 
                           registers_25_26_port, B2 => n4934, ZN => n1455);
   U1372 : AOI22_X1 port map( A1 => registers_12_25_port, A2 => n4961, B1 => 
                           registers_30_25_port, B2 => n4958, ZN => n1416);
   U1373 : AOI22_X1 port map( A1 => registers_20_25_port, A2 => n4949, B1 => 
                           registers_21_25_port, B2 => n4946, ZN => n1419);
   U1374 : AOI22_X1 port map( A1 => registers_24_25_port, A2 => n4937, B1 => 
                           registers_25_25_port, B2 => n4934, ZN => n1422);
   U1375 : AOI22_X1 port map( A1 => registers_12_24_port, A2 => n4961, B1 => 
                           registers_30_24_port, B2 => n4958, ZN => n1383);
   U1376 : AOI22_X1 port map( A1 => registers_20_24_port, A2 => n4949, B1 => 
                           registers_21_24_port, B2 => n4946, ZN => n1386);
   U1377 : AOI22_X1 port map( A1 => registers_24_24_port, A2 => n4937, B1 => 
                           registers_25_24_port, B2 => n4934, ZN => n1389);
   U1378 : AOI22_X1 port map( A1 => registers_12_23_port, A2 => n4961, B1 => 
                           registers_30_23_port, B2 => n4958, ZN => n1350);
   U1379 : AOI22_X1 port map( A1 => registers_20_23_port, A2 => n4949, B1 => 
                           registers_21_23_port, B2 => n4946, ZN => n1353);
   U1380 : AOI22_X1 port map( A1 => registers_24_23_port, A2 => n4937, B1 => 
                           registers_25_23_port, B2 => n4934, ZN => n1356);
   U1381 : AOI22_X1 port map( A1 => registers_12_22_port, A2 => n4961, B1 => 
                           registers_30_22_port, B2 => n4958, ZN => n1317);
   U1382 : AOI22_X1 port map( A1 => registers_20_22_port, A2 => n4949, B1 => 
                           registers_21_22_port, B2 => n4946, ZN => n1320);
   U1383 : AOI22_X1 port map( A1 => registers_24_22_port, A2 => n4937, B1 => 
                           registers_25_22_port, B2 => n4934, ZN => n1323);
   U1384 : AOI22_X1 port map( A1 => registers_12_21_port, A2 => n4961, B1 => 
                           registers_30_21_port, B2 => n4958, ZN => n1284);
   U1385 : AOI22_X1 port map( A1 => registers_20_21_port, A2 => n4949, B1 => 
                           registers_21_21_port, B2 => n4946, ZN => n1287);
   U1386 : AOI22_X1 port map( A1 => registers_24_21_port, A2 => n4937, B1 => 
                           registers_25_21_port, B2 => n4934, ZN => n1290);
   U1387 : AOI22_X1 port map( A1 => registers_12_20_port, A2 => n4961, B1 => 
                           registers_30_20_port, B2 => n4958, ZN => n1251);
   U1388 : AOI22_X1 port map( A1 => registers_20_20_port, A2 => n4949, B1 => 
                           registers_21_20_port, B2 => n4946, ZN => n1254);
   U1389 : AOI22_X1 port map( A1 => registers_24_20_port, A2 => n4937, B1 => 
                           registers_25_20_port, B2 => n4934, ZN => n1257);
   U1390 : AOI22_X1 port map( A1 => registers_12_19_port, A2 => n4962, B1 => 
                           registers_30_19_port, B2 => n4959, ZN => n1218);
   U1391 : AOI22_X1 port map( A1 => registers_20_19_port, A2 => n4950, B1 => 
                           registers_21_19_port, B2 => n4947, ZN => n1221);
   U1392 : AOI22_X1 port map( A1 => registers_24_19_port, A2 => n4938, B1 => 
                           registers_25_19_port, B2 => n4935, ZN => n1224);
   U1393 : AOI22_X1 port map( A1 => registers_12_18_port, A2 => n4962, B1 => 
                           registers_30_18_port, B2 => n4959, ZN => n1185);
   U1394 : AOI22_X1 port map( A1 => registers_20_18_port, A2 => n4950, B1 => 
                           registers_21_18_port, B2 => n4947, ZN => n1188);
   U1395 : AOI22_X1 port map( A1 => registers_24_18_port, A2 => n4938, B1 => 
                           registers_25_18_port, B2 => n4935, ZN => n1191);
   U1396 : AOI22_X1 port map( A1 => registers_12_17_port, A2 => n4962, B1 => 
                           registers_30_17_port, B2 => n4959, ZN => n1152);
   U1397 : AOI22_X1 port map( A1 => registers_20_17_port, A2 => n4950, B1 => 
                           registers_21_17_port, B2 => n4947, ZN => n1155);
   U1398 : AOI22_X1 port map( A1 => registers_24_17_port, A2 => n4938, B1 => 
                           registers_25_17_port, B2 => n4935, ZN => n1158);
   U1399 : AOI22_X1 port map( A1 => registers_12_16_port, A2 => n4962, B1 => 
                           registers_30_16_port, B2 => n4959, ZN => n1119);
   U1400 : AOI22_X1 port map( A1 => registers_20_16_port, A2 => n4950, B1 => 
                           registers_21_16_port, B2 => n4947, ZN => n1122);
   U1401 : AOI22_X1 port map( A1 => registers_24_16_port, A2 => n4938, B1 => 
                           registers_25_16_port, B2 => n4935, ZN => n1125);
   U1402 : INV_X1 port map( A => address_port_a(4), ZN => n1637);
   U1403 : INV_X1 port map( A => address_port_b(0), ZN => n2302);
   U1404 : INV_X1 port map( A => address_port_a(0), ZN => n1642);
   U1405 : INV_X1 port map( A => address_port_a(3), ZN => n1641);
   U1406 : INV_X1 port map( A => address_port_b(4), ZN => n2299);
   U1407 : INV_X1 port map( A => address_port_b(3), ZN => n2301);
   U1408 : NAND4_X1 port map( A1 => n809, A2 => n810, A3 => n811, A4 => n812, 
                           ZN => n1836);
   U1409 : AOI211_X1 port map( C1 => registers_15_7_port, C2 => n4933, A => 
                           n829, B => n830, ZN => n811);
   U1410 : AOI221_X1 port map( B1 => registers_29_7_port, B2 => n4900, C1 => 
                           registers_10_7_port, C2 => n4897, A => n839, ZN => 
                           n809);
   U1411 : AOI221_X1 port map( B1 => registers_27_7_port, B2 => n4912, C1 => 
                           registers_7_7_port, C2 => n4909, A => n836, ZN => 
                           n810);
   U1412 : NAND4_X1 port map( A1 => n776, A2 => n777, A3 => n778, A4 => n779, 
                           ZN => n1837);
   U1413 : AOI211_X1 port map( C1 => registers_15_6_port, C2 => n4933, A => 
                           n796, B => n797, ZN => n778);
   U1414 : AOI221_X1 port map( B1 => registers_29_6_port, B2 => n4900, C1 => 
                           registers_10_6_port, C2 => n4897, A => n806, ZN => 
                           n776);
   U1415 : AOI221_X1 port map( B1 => registers_27_6_port, B2 => n4912, C1 => 
                           registers_7_6_port, C2 => n4909, A => n803, ZN => 
                           n777);
   U1416 : NAND4_X1 port map( A1 => n743, A2 => n744, A3 => n745, A4 => n746, 
                           ZN => n1838);
   U1417 : AOI211_X1 port map( C1 => registers_15_5_port, C2 => n4933, A => 
                           n763, B => n764, ZN => n745);
   U1418 : AOI221_X1 port map( B1 => registers_29_5_port, B2 => n4900, C1 => 
                           registers_10_5_port, C2 => n4897, A => n773, ZN => 
                           n743);
   U1419 : AOI221_X1 port map( B1 => registers_27_5_port, B2 => n4912, C1 => 
                           registers_7_5_port, C2 => n4909, A => n770, ZN => 
                           n744);
   U1420 : NAND4_X1 port map( A1 => n710, A2 => n711, A3 => n712, A4 => n713, 
                           ZN => n1839);
   U1421 : AOI211_X1 port map( C1 => registers_15_4_port, C2 => n4933, A => 
                           n730, B => n731, ZN => n712);
   U1422 : AOI221_X1 port map( B1 => registers_29_4_port, B2 => n4900, C1 => 
                           registers_10_4_port, C2 => n4897, A => n740, ZN => 
                           n710);
   U1423 : AOI221_X1 port map( B1 => registers_27_4_port, B2 => n4912, C1 => 
                           registers_7_4_port, C2 => n4909, A => n737, ZN => 
                           n711);
   U1424 : NAND4_X1 port map( A1 => n677, A2 => n678, A3 => n679, A4 => n680, 
                           ZN => n1840);
   U1425 : AOI211_X1 port map( C1 => registers_15_3_port, C2 => n4933, A => 
                           n697, B => n698, ZN => n679);
   U1426 : AOI221_X1 port map( B1 => registers_29_3_port, B2 => n4900, C1 => 
                           registers_10_3_port, C2 => n4897, A => n707, ZN => 
                           n677);
   U1427 : AOI221_X1 port map( B1 => registers_27_3_port, B2 => n4912, C1 => 
                           registers_7_3_port, C2 => n4909, A => n704, ZN => 
                           n678);
   U1428 : NAND4_X1 port map( A1 => n644, A2 => n645, A3 => n646, A4 => n647, 
                           ZN => n1841);
   U1429 : AOI211_X1 port map( C1 => registers_15_2_port, C2 => n4933, A => 
                           n664, B => n665, ZN => n646);
   U1430 : AOI221_X1 port map( B1 => registers_29_2_port, B2 => n4900, C1 => 
                           registers_10_2_port, C2 => n4897, A => n674, ZN => 
                           n644);
   U1431 : AOI221_X1 port map( B1 => registers_27_2_port, B2 => n4912, C1 => 
                           registers_7_2_port, C2 => n4909, A => n671, ZN => 
                           n645);
   U1432 : NAND4_X1 port map( A1 => n611, A2 => n612, A3 => n613, A4 => n614, 
                           ZN => n1842);
   U1433 : AOI211_X1 port map( C1 => registers_15_1_port, C2 => n4933, A => 
                           n631, B => n632, ZN => n613);
   U1434 : AOI221_X1 port map( B1 => registers_29_1_port, B2 => n4900, C1 => 
                           registers_10_1_port, C2 => n4897, A => n641, ZN => 
                           n611);
   U1435 : AOI221_X1 port map( B1 => registers_27_1_port, B2 => n4912, C1 => 
                           registers_7_1_port, C2 => n4909, A => n638, ZN => 
                           n612);
   U1436 : NAND4_X1 port map( A1 => n547, A2 => n548, A3 => n549, A4 => n550, 
                           ZN => n1843);
   U1437 : AOI211_X1 port map( C1 => registers_15_0_port, C2 => n4933, A => 
                           n584, B => n585, ZN => n549);
   U1438 : AOI221_X1 port map( B1 => registers_29_0_port, B2 => n4900, C1 => 
                           registers_10_0_port, C2 => n4897, A => n606, ZN => 
                           n547);
   U1439 : AOI221_X1 port map( B1 => registers_27_0_port, B2 => n4912, C1 => 
                           registers_7_0_port, C2 => n4909, A => n599, ZN => 
                           n548);
   U1440 : NAND4_X1 port map( A1 => n2001, A2 => n2002, A3 => n2003, A4 => 
                           n2004, ZN => n1794);
   U1441 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_15_port, A => 
                           n2013, B => n2014, ZN => n2003);
   U1442 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_15_port, C1 => 
                           n4803, C2 => registers_10_15_port, A => n2017, ZN =>
                           n2001);
   U1443 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_15_port, C1 => 
                           n4815, C2 => registers_7_15_port, A => n2016, ZN => 
                           n2002);
   U1444 : NAND4_X1 port map( A1 => n1984, A2 => n1985, A3 => n1986, A4 => 
                           n1987, ZN => n1795);
   U1445 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_14_port, A => 
                           n1996, B => n1997, ZN => n1986);
   U1446 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_14_port, C1 => 
                           n4803, C2 => registers_10_14_port, A => n2000, ZN =>
                           n1984);
   U1447 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_14_port, C1 => 
                           n4815, C2 => registers_7_14_port, A => n1999, ZN => 
                           n1985);
   U1448 : NAND4_X1 port map( A1 => n1967, A2 => n1968, A3 => n1969, A4 => 
                           n1970, ZN => n1796);
   U1449 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_13_port, A => 
                           n1979, B => n1980, ZN => n1969);
   U1450 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_13_port, C1 => 
                           n4803, C2 => registers_10_13_port, A => n1983, ZN =>
                           n1967);
   U1451 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_13_port, C1 => 
                           n4815, C2 => registers_7_13_port, A => n1982, ZN => 
                           n1968);
   U1452 : NAND4_X1 port map( A1 => n1950, A2 => n1951, A3 => n1952, A4 => 
                           n1953, ZN => n1797);
   U1453 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_12_port, A => 
                           n1962, B => n1963, ZN => n1952);
   U1454 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_12_port, C1 => 
                           n4803, C2 => registers_10_12_port, A => n1966, ZN =>
                           n1950);
   U1455 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_12_port, C1 => 
                           n4815, C2 => registers_7_12_port, A => n1965, ZN => 
                           n1951);
   U1456 : NAND4_X1 port map( A1 => n1933, A2 => n1934, A3 => n1935, A4 => 
                           n1936, ZN => n1798);
   U1457 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_11_port, A => 
                           n1945, B => n1946, ZN => n1935);
   U1458 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_11_port, C1 => 
                           n4803, C2 => registers_10_11_port, A => n1949, ZN =>
                           n1933);
   U1459 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_11_port, C1 => 
                           n4815, C2 => registers_7_11_port, A => n1948, ZN => 
                           n1934);
   U1460 : NAND4_X1 port map( A1 => n1916, A2 => n1917, A3 => n1918, A4 => 
                           n1919, ZN => n1799);
   U1461 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_10_port, A => 
                           n1928, B => n1929, ZN => n1918);
   U1462 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_10_port, C1 => 
                           n4803, C2 => registers_10_10_port, A => n1932, ZN =>
                           n1916);
   U1463 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_10_port, C1 => 
                           n4815, C2 => registers_7_10_port, A => n1931, ZN => 
                           n1917);
   U1464 : NAND4_X1 port map( A1 => n1899, A2 => n1900, A3 => n1901, A4 => 
                           n1902, ZN => n1800);
   U1465 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_9_port, A => 
                           n1911, B => n1912, ZN => n1901);
   U1466 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_9_port, C1 => 
                           n4803, C2 => registers_10_9_port, A => n1915, ZN => 
                           n1899);
   U1467 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_9_port, C1 => 
                           n4815, C2 => registers_7_9_port, A => n1914, ZN => 
                           n1900);
   U1468 : NAND4_X1 port map( A1 => n1882, A2 => n1883, A3 => n1884, A4 => 
                           n1885, ZN => n1802);
   U1469 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_8_port, A => 
                           n1894, B => n1895, ZN => n1884);
   U1470 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_8_port, C1 => 
                           n4803, C2 => registers_10_8_port, A => n1898, ZN => 
                           n1882);
   U1471 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_8_port, C1 => 
                           n4815, C2 => registers_7_8_port, A => n1897, ZN => 
                           n1883);
   U1472 : NAND4_X1 port map( A1 => n1073, A2 => n1074, A3 => n1075, A4 => 
                           n1076, ZN => n1827);
   U1473 : AOI211_X1 port map( C1 => registers_15_15_port, C2 => n4932, A => 
                           n1093, B => n1094, ZN => n1075);
   U1474 : AOI221_X1 port map( B1 => registers_29_15_port, B2 => n4899, C1 => 
                           registers_10_15_port, C2 => n4896, A => n1103, ZN =>
                           n1073);
   U1475 : AOI221_X1 port map( B1 => registers_27_15_port, B2 => n4911, C1 => 
                           registers_7_15_port, C2 => n4908, A => n1100, ZN => 
                           n1074);
   U1476 : NAND4_X1 port map( A1 => n1040, A2 => n1041, A3 => n1042, A4 => 
                           n1043, ZN => n1828);
   U1477 : AOI211_X1 port map( C1 => registers_15_14_port, C2 => n4932, A => 
                           n1060, B => n1061, ZN => n1042);
   U1478 : AOI221_X1 port map( B1 => registers_29_14_port, B2 => n4899, C1 => 
                           registers_10_14_port, C2 => n4896, A => n1070, ZN =>
                           n1040);
   U1479 : AOI221_X1 port map( B1 => registers_27_14_port, B2 => n4911, C1 => 
                           registers_7_14_port, C2 => n4908, A => n1067, ZN => 
                           n1041);
   U1480 : NAND4_X1 port map( A1 => n1007, A2 => n1008, A3 => n1009, A4 => 
                           n1010, ZN => n1829);
   U1481 : AOI211_X1 port map( C1 => registers_15_13_port, C2 => n4932, A => 
                           n1027, B => n1028, ZN => n1009);
   U1482 : AOI221_X1 port map( B1 => registers_29_13_port, B2 => n4899, C1 => 
                           registers_10_13_port, C2 => n4896, A => n1037, ZN =>
                           n1007);
   U1483 : AOI221_X1 port map( B1 => registers_27_13_port, B2 => n4911, C1 => 
                           registers_7_13_port, C2 => n4908, A => n1034, ZN => 
                           n1008);
   U1484 : NAND4_X1 port map( A1 => n974, A2 => n975, A3 => n976, A4 => n977, 
                           ZN => n1830);
   U1485 : AOI211_X1 port map( C1 => registers_15_12_port, C2 => n4932, A => 
                           n994, B => n995, ZN => n976);
   U1486 : AOI221_X1 port map( B1 => registers_29_12_port, B2 => n4899, C1 => 
                           registers_10_12_port, C2 => n4896, A => n1004, ZN =>
                           n974);
   U1487 : AOI221_X1 port map( B1 => registers_27_12_port, B2 => n4911, C1 => 
                           registers_7_12_port, C2 => n4908, A => n1001, ZN => 
                           n975);
   U1488 : NAND4_X1 port map( A1 => n941, A2 => n942, A3 => n943, A4 => n944, 
                           ZN => n1831);
   U1489 : AOI211_X1 port map( C1 => registers_15_11_port, C2 => n4932, A => 
                           n961, B => n962, ZN => n943);
   U1490 : AOI221_X1 port map( B1 => registers_29_11_port, B2 => n4899, C1 => 
                           registers_10_11_port, C2 => n4896, A => n971, ZN => 
                           n941);
   U1491 : AOI221_X1 port map( B1 => registers_27_11_port, B2 => n4911, C1 => 
                           registers_7_11_port, C2 => n4908, A => n968, ZN => 
                           n942);
   U1492 : NAND4_X1 port map( A1 => n908, A2 => n909, A3 => n910, A4 => n911, 
                           ZN => n1832);
   U1493 : AOI211_X1 port map( C1 => registers_15_10_port, C2 => n4932, A => 
                           n928, B => n929, ZN => n910);
   U1494 : AOI221_X1 port map( B1 => registers_29_10_port, B2 => n4899, C1 => 
                           registers_10_10_port, C2 => n4896, A => n938, ZN => 
                           n908);
   U1495 : AOI221_X1 port map( B1 => registers_27_10_port, B2 => n4911, C1 => 
                           registers_7_10_port, C2 => n4908, A => n935, ZN => 
                           n909);
   U1496 : NAND4_X1 port map( A1 => n875, A2 => n876, A3 => n877, A4 => n878, 
                           ZN => n1833);
   U1497 : AOI211_X1 port map( C1 => registers_15_9_port, C2 => n4932, A => 
                           n895, B => n896, ZN => n877);
   U1498 : AOI221_X1 port map( B1 => registers_29_9_port, B2 => n4899, C1 => 
                           registers_10_9_port, C2 => n4896, A => n905, ZN => 
                           n875);
   U1499 : AOI221_X1 port map( B1 => registers_27_9_port, B2 => n4911, C1 => 
                           registers_7_9_port, C2 => n4908, A => n902, ZN => 
                           n876);
   U1500 : NAND4_X1 port map( A1 => n842, A2 => n843, A3 => n844, A4 => n845, 
                           ZN => n1835);
   U1501 : AOI211_X1 port map( C1 => registers_15_8_port, C2 => n4932, A => 
                           n862, B => n863, ZN => n844);
   U1502 : AOI221_X1 port map( B1 => registers_29_8_port, B2 => n4899, C1 => 
                           registers_10_8_port, C2 => n4896, A => n872, ZN => 
                           n842);
   U1503 : AOI221_X1 port map( B1 => registers_27_8_port, B2 => n4911, C1 => 
                           registers_7_8_port, C2 => n4908, A => n869, ZN => 
                           n843);
   U1504 : NAND4_X1 port map( A1 => n1865, A2 => n1866, A3 => n1867, A4 => 
                           n1868, ZN => n1803);
   U1505 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_7_port, A => 
                           n1877, B => n1878, ZN => n1867);
   U1506 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_7_port, C1 => 
                           n4804, C2 => registers_10_7_port, A => n1881, ZN => 
                           n1865);
   U1507 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_7_port, C1 => 
                           n4816, C2 => registers_7_7_port, A => n1880, ZN => 
                           n1866);
   U1508 : NAND4_X1 port map( A1 => n1848, A2 => n1849, A3 => n1850, A4 => 
                           n1851, ZN => n1804);
   U1509 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_6_port, A => 
                           n1860, B => n1861, ZN => n1850);
   U1510 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_6_port, C1 => 
                           n4804, C2 => registers_10_6_port, A => n1864, ZN => 
                           n1848);
   U1511 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_6_port, C1 => 
                           n4816, C2 => registers_7_6_port, A => n1863, ZN => 
                           n1849);
   U1512 : NAND4_X1 port map( A1 => n1767, A2 => n1768, A3 => n1769, A4 => 
                           n1770, ZN => n1805);
   U1513 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_5_port, A => 
                           n1834, B => n1844, ZN => n1769);
   U1514 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_5_port, C1 => 
                           n4804, C2 => registers_10_5_port, A => n1847, ZN => 
                           n1767);
   U1515 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_5_port, C1 => 
                           n4816, C2 => registers_7_5_port, A => n1846, ZN => 
                           n1768);
   U1516 : NAND4_X1 port map( A1 => n1750, A2 => n1751, A3 => n1752, A4 => 
                           n1753, ZN => n1806);
   U1517 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_4_port, A => 
                           n1762, B => n1763, ZN => n1752);
   U1518 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_4_port, C1 => 
                           n4804, C2 => registers_10_4_port, A => n1766, ZN => 
                           n1750);
   U1519 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_4_port, C1 => 
                           n4816, C2 => registers_7_4_port, A => n1765, ZN => 
                           n1751);
   U1520 : NAND4_X1 port map( A1 => n1733, A2 => n1734, A3 => n1735, A4 => 
                           n1736, ZN => n1807);
   U1521 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_3_port, A => 
                           n1745, B => n1746, ZN => n1735);
   U1522 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_3_port, C1 => 
                           n4804, C2 => registers_10_3_port, A => n1749, ZN => 
                           n1733);
   U1523 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_3_port, C1 => 
                           n4816, C2 => registers_7_3_port, A => n1748, ZN => 
                           n1734);
   U1524 : NAND4_X1 port map( A1 => n1716, A2 => n1717, A3 => n1718, A4 => 
                           n1719, ZN => n1808);
   U1525 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_2_port, A => 
                           n1728, B => n1729, ZN => n1718);
   U1526 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_2_port, C1 => 
                           n4804, C2 => registers_10_2_port, A => n1732, ZN => 
                           n1716);
   U1527 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_2_port, C1 => 
                           n4816, C2 => registers_7_2_port, A => n1731, ZN => 
                           n1717);
   U1528 : NAND4_X1 port map( A1 => n1699, A2 => n1700, A3 => n1701, A4 => 
                           n1702, ZN => n1809);
   U1529 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_1_port, A => 
                           n1711, B => n1712, ZN => n1701);
   U1530 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_1_port, C1 => 
                           n4804, C2 => registers_10_1_port, A => n1715, ZN => 
                           n1699);
   U1531 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_1_port, C1 => 
                           n4816, C2 => registers_7_1_port, A => n1714, ZN => 
                           n1700);
   U1532 : NAND4_X1 port map( A1 => n1651, A2 => n1652, A3 => n1653, A4 => 
                           n1654, ZN => n1810);
   U1533 : AOI211_X1 port map( C1 => n4840, C2 => registers_15_0_port, A => 
                           n1680, B => n1681, ZN => n1653);
   U1534 : AOI221_X1 port map( B1 => n4807, B2 => registers_29_0_port, C1 => 
                           n4804, C2 => registers_10_0_port, A => n1696, ZN => 
                           n1651);
   U1535 : AOI221_X1 port map( B1 => n4819, B2 => registers_27_0_port, C1 => 
                           n4816, C2 => registers_7_0_port, A => n1691, ZN => 
                           n1652);
   U1536 : NAND4_X1 port map( A1 => n2273, A2 => n2274, A3 => n2275, A4 => 
                           n2276, ZN => n1778);
   U1537 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_31_port, A => 
                           n2297, B => n2298, ZN => n2275);
   U1538 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_31_port, C1 => 
                           n4802, C2 => registers_10_31_port, A => n2304, ZN =>
                           n2273);
   U1539 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_31_port, C1 => 
                           n4814, C2 => registers_7_31_port, A => n2303, ZN => 
                           n2274);
   U1540 : NAND4_X1 port map( A1 => n2256, A2 => n2257, A3 => n2258, A4 => 
                           n2259, ZN => n1779);
   U1541 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_30_port, A => 
                           n2268, B => n2269, ZN => n2258);
   U1542 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_30_port, C1 => 
                           n4802, C2 => registers_10_30_port, A => n2272, ZN =>
                           n2256);
   U1543 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_30_port, C1 => 
                           n4814, C2 => registers_7_30_port, A => n2271, ZN => 
                           n2257);
   U1544 : NAND4_X1 port map( A1 => n2239, A2 => n2240, A3 => n2241, A4 => 
                           n2242, ZN => n1780);
   U1545 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_29_port, A => 
                           n2251, B => n2252, ZN => n2241);
   U1546 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_29_port, C1 => 
                           n4802, C2 => registers_10_29_port, A => n2255, ZN =>
                           n2239);
   U1547 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_29_port, C1 => 
                           n4814, C2 => registers_7_29_port, A => n2254, ZN => 
                           n2240);
   U1548 : NAND4_X1 port map( A1 => n2222, A2 => n2223, A3 => n2224, A4 => 
                           n2225, ZN => n1781);
   U1549 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_28_port, A => 
                           n2234, B => n2235, ZN => n2224);
   U1550 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_28_port, C1 => 
                           n4802, C2 => registers_10_28_port, A => n2238, ZN =>
                           n2222);
   U1551 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_28_port, C1 => 
                           n4814, C2 => registers_7_28_port, A => n2237, ZN => 
                           n2223);
   U1552 : NAND4_X1 port map( A1 => n2205, A2 => n2206, A3 => n2207, A4 => 
                           n2208, ZN => n1782);
   U1553 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_27_port, A => 
                           n2217, B => n2218, ZN => n2207);
   U1554 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_27_port, C1 => 
                           n4802, C2 => registers_10_27_port, A => n2221, ZN =>
                           n2205);
   U1555 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_27_port, C1 => 
                           n4814, C2 => registers_7_27_port, A => n2220, ZN => 
                           n2206);
   U1556 : NAND4_X1 port map( A1 => n2188, A2 => n2189, A3 => n2190, A4 => 
                           n2191, ZN => n1783);
   U1557 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_26_port, A => 
                           n2200, B => n2201, ZN => n2190);
   U1558 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_26_port, C1 => 
                           n4802, C2 => registers_10_26_port, A => n2204, ZN =>
                           n2188);
   U1559 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_26_port, C1 => 
                           n4814, C2 => registers_7_26_port, A => n2203, ZN => 
                           n2189);
   U1560 : NAND4_X1 port map( A1 => n2171, A2 => n2172, A3 => n2173, A4 => 
                           n2174, ZN => n1784);
   U1561 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_25_port, A => 
                           n2183, B => n2184, ZN => n2173);
   U1562 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_25_port, C1 => 
                           n4802, C2 => registers_10_25_port, A => n2187, ZN =>
                           n2171);
   U1563 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_25_port, C1 => 
                           n4814, C2 => registers_7_25_port, A => n2186, ZN => 
                           n2172);
   U1564 : NAND4_X1 port map( A1 => n2154, A2 => n2155, A3 => n2156, A4 => 
                           n2157, ZN => n1785);
   U1565 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_24_port, A => 
                           n2166, B => n2167, ZN => n2156);
   U1566 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_24_port, C1 => 
                           n4802, C2 => registers_10_24_port, A => n2170, ZN =>
                           n2154);
   U1567 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_24_port, C1 => 
                           n4814, C2 => registers_7_24_port, A => n2169, ZN => 
                           n2155);
   U1568 : NAND4_X1 port map( A1 => n2137, A2 => n2138, A3 => n2139, A4 => 
                           n2140, ZN => n1786);
   U1569 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_23_port, A => 
                           n2149, B => n2150, ZN => n2139);
   U1570 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_23_port, C1 => 
                           n4802, C2 => registers_10_23_port, A => n2153, ZN =>
                           n2137);
   U1571 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_23_port, C1 => 
                           n4814, C2 => registers_7_23_port, A => n2152, ZN => 
                           n2138);
   U1572 : NAND4_X1 port map( A1 => n2120, A2 => n2121, A3 => n2122, A4 => 
                           n2123, ZN => n1787);
   U1573 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_22_port, A => 
                           n2132, B => n2133, ZN => n2122);
   U1574 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_22_port, C1 => 
                           n4802, C2 => registers_10_22_port, A => n2136, ZN =>
                           n2120);
   U1575 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_22_port, C1 => 
                           n4814, C2 => registers_7_22_port, A => n2135, ZN => 
                           n2121);
   U1576 : NAND4_X1 port map( A1 => n2103, A2 => n2104, A3 => n2105, A4 => 
                           n2106, ZN => n1788);
   U1577 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_21_port, A => 
                           n2115, B => n2116, ZN => n2105);
   U1578 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_21_port, C1 => 
                           n4802, C2 => registers_10_21_port, A => n2119, ZN =>
                           n2103);
   U1579 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_21_port, C1 => 
                           n4814, C2 => registers_7_21_port, A => n2118, ZN => 
                           n2104);
   U1580 : NAND4_X1 port map( A1 => n2086, A2 => n2087, A3 => n2088, A4 => 
                           n2089, ZN => n1789);
   U1581 : AOI211_X1 port map( C1 => n4838, C2 => registers_15_20_port, A => 
                           n2098, B => n2099, ZN => n2088);
   U1582 : AOI221_X1 port map( B1 => n4805, B2 => registers_29_20_port, C1 => 
                           n4802, C2 => registers_10_20_port, A => n2102, ZN =>
                           n2086);
   U1583 : AOI221_X1 port map( B1 => n4817, B2 => registers_27_20_port, C1 => 
                           n4814, C2 => registers_7_20_port, A => n2101, ZN => 
                           n2087);
   U1584 : NAND4_X1 port map( A1 => n2069, A2 => n2070, A3 => n2071, A4 => 
                           n2072, ZN => n1790);
   U1585 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_19_port, A => 
                           n2081, B => n2082, ZN => n2071);
   U1586 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_19_port, C1 => 
                           n4803, C2 => registers_10_19_port, A => n2085, ZN =>
                           n2069);
   U1587 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_19_port, C1 => 
                           n4815, C2 => registers_7_19_port, A => n2084, ZN => 
                           n2070);
   U1588 : NAND4_X1 port map( A1 => n2052, A2 => n2053, A3 => n2054, A4 => 
                           n2055, ZN => n1791);
   U1589 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_18_port, A => 
                           n2064, B => n2065, ZN => n2054);
   U1590 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_18_port, C1 => 
                           n4803, C2 => registers_10_18_port, A => n2068, ZN =>
                           n2052);
   U1591 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_18_port, C1 => 
                           n4815, C2 => registers_7_18_port, A => n2067, ZN => 
                           n2053);
   U1592 : NAND4_X1 port map( A1 => n2035, A2 => n2036, A3 => n2037, A4 => 
                           n2038, ZN => n1792);
   U1593 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_17_port, A => 
                           n2047, B => n2048, ZN => n2037);
   U1594 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_17_port, C1 => 
                           n4803, C2 => registers_10_17_port, A => n2051, ZN =>
                           n2035);
   U1595 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_17_port, C1 => 
                           n4815, C2 => registers_7_17_port, A => n2050, ZN => 
                           n2036);
   U1596 : NAND4_X1 port map( A1 => n2018, A2 => n2019, A3 => n2020, A4 => 
                           n2021, ZN => n1793);
   U1597 : AOI211_X1 port map( C1 => n4839, C2 => registers_15_16_port, A => 
                           n2030, B => n2031, ZN => n2020);
   U1598 : AOI221_X1 port map( B1 => n4806, B2 => registers_29_16_port, C1 => 
                           n4803, C2 => registers_10_16_port, A => n2034, ZN =>
                           n2018);
   U1599 : AOI221_X1 port map( B1 => n4818, B2 => registers_27_16_port, C1 => 
                           n4815, C2 => registers_7_16_port, A => n2033, ZN => 
                           n2019);
   U1600 : NAND4_X1 port map( A1 => n1601, A2 => n1602, A3 => n1603, A4 => 
                           n1604, ZN => n1811);
   U1601 : AOI211_X1 port map( C1 => registers_15_31_port, C2 => n4931, A => 
                           n1633, B => n1634, ZN => n1603);
   U1602 : AOI221_X1 port map( B1 => registers_29_31_port, B2 => n4898, C1 => 
                           registers_10_31_port, C2 => n4895, A => n1646, ZN =>
                           n1601);
   U1603 : AOI221_X1 port map( B1 => registers_27_31_port, B2 => n4910, C1 => 
                           registers_7_31_port, C2 => n4907, A => n1643, ZN => 
                           n1602);
   U1604 : NAND4_X1 port map( A1 => n1568, A2 => n1569, A3 => n1570, A4 => 
                           n1571, ZN => n1812);
   U1605 : AOI211_X1 port map( C1 => registers_15_30_port, C2 => n4931, A => 
                           n1588, B => n1589, ZN => n1570);
   U1606 : AOI221_X1 port map( B1 => registers_29_30_port, B2 => n4898, C1 => 
                           registers_10_30_port, C2 => n4895, A => n1598, ZN =>
                           n1568);
   U1607 : AOI221_X1 port map( B1 => registers_27_30_port, B2 => n4910, C1 => 
                           registers_7_30_port, C2 => n4907, A => n1595, ZN => 
                           n1569);
   U1608 : NAND4_X1 port map( A1 => n1535, A2 => n1536, A3 => n1537, A4 => 
                           n1538, ZN => n1813);
   U1609 : AOI211_X1 port map( C1 => registers_15_29_port, C2 => n4931, A => 
                           n1555, B => n1556, ZN => n1537);
   U1610 : AOI221_X1 port map( B1 => registers_29_29_port, B2 => n4898, C1 => 
                           registers_10_29_port, C2 => n4895, A => n1565, ZN =>
                           n1535);
   U1611 : AOI221_X1 port map( B1 => registers_27_29_port, B2 => n4910, C1 => 
                           registers_7_29_port, C2 => n4907, A => n1562, ZN => 
                           n1536);
   U1612 : NAND4_X1 port map( A1 => n1502, A2 => n1503, A3 => n1504, A4 => 
                           n1505, ZN => n1814);
   U1613 : AOI211_X1 port map( C1 => registers_15_28_port, C2 => n4931, A => 
                           n1522, B => n1523, ZN => n1504);
   U1614 : AOI221_X1 port map( B1 => registers_29_28_port, B2 => n4898, C1 => 
                           registers_10_28_port, C2 => n4895, A => n1532, ZN =>
                           n1502);
   U1615 : AOI221_X1 port map( B1 => registers_27_28_port, B2 => n4910, C1 => 
                           registers_7_28_port, C2 => n4907, A => n1529, ZN => 
                           n1503);
   U1616 : NAND4_X1 port map( A1 => n1469, A2 => n1470, A3 => n1471, A4 => 
                           n1472, ZN => n1815);
   U1617 : AOI211_X1 port map( C1 => registers_15_27_port, C2 => n4931, A => 
                           n1489, B => n1490, ZN => n1471);
   U1618 : AOI221_X1 port map( B1 => registers_29_27_port, B2 => n4898, C1 => 
                           registers_10_27_port, C2 => n4895, A => n1499, ZN =>
                           n1469);
   U1619 : AOI221_X1 port map( B1 => registers_27_27_port, B2 => n4910, C1 => 
                           registers_7_27_port, C2 => n4907, A => n1496, ZN => 
                           n1470);
   U1620 : NAND4_X1 port map( A1 => n1436, A2 => n1437, A3 => n1438, A4 => 
                           n1439, ZN => n1816);
   U1621 : AOI211_X1 port map( C1 => registers_15_26_port, C2 => n4931, A => 
                           n1456, B => n1457, ZN => n1438);
   U1622 : AOI221_X1 port map( B1 => registers_29_26_port, B2 => n4898, C1 => 
                           registers_10_26_port, C2 => n4895, A => n1466, ZN =>
                           n1436);
   U1623 : AOI221_X1 port map( B1 => registers_27_26_port, B2 => n4910, C1 => 
                           registers_7_26_port, C2 => n4907, A => n1463, ZN => 
                           n1437);
   U1624 : NAND4_X1 port map( A1 => n1403, A2 => n1404, A3 => n1405, A4 => 
                           n1406, ZN => n1817);
   U1625 : AOI211_X1 port map( C1 => registers_15_25_port, C2 => n4931, A => 
                           n1423, B => n1424, ZN => n1405);
   U1626 : AOI221_X1 port map( B1 => registers_29_25_port, B2 => n4898, C1 => 
                           registers_10_25_port, C2 => n4895, A => n1433, ZN =>
                           n1403);
   U1627 : AOI221_X1 port map( B1 => registers_27_25_port, B2 => n4910, C1 => 
                           registers_7_25_port, C2 => n4907, A => n1430, ZN => 
                           n1404);
   U1628 : NAND4_X1 port map( A1 => n1370, A2 => n1371, A3 => n1372, A4 => 
                           n1373, ZN => n1818);
   U1629 : AOI211_X1 port map( C1 => registers_15_24_port, C2 => n4931, A => 
                           n1390, B => n1391, ZN => n1372);
   U1630 : AOI221_X1 port map( B1 => registers_29_24_port, B2 => n4898, C1 => 
                           registers_10_24_port, C2 => n4895, A => n1400, ZN =>
                           n1370);
   U1631 : AOI221_X1 port map( B1 => registers_27_24_port, B2 => n4910, C1 => 
                           registers_7_24_port, C2 => n4907, A => n1397, ZN => 
                           n1371);
   U1632 : NAND4_X1 port map( A1 => n1337, A2 => n1338, A3 => n1339, A4 => 
                           n1340, ZN => n1819);
   U1633 : AOI211_X1 port map( C1 => registers_15_23_port, C2 => n4931, A => 
                           n1357, B => n1358, ZN => n1339);
   U1634 : AOI221_X1 port map( B1 => registers_29_23_port, B2 => n4898, C1 => 
                           registers_10_23_port, C2 => n4895, A => n1367, ZN =>
                           n1337);
   U1635 : AOI221_X1 port map( B1 => registers_27_23_port, B2 => n4910, C1 => 
                           registers_7_23_port, C2 => n4907, A => n1364, ZN => 
                           n1338);
   U1636 : NAND4_X1 port map( A1 => n1304, A2 => n1305, A3 => n1306, A4 => 
                           n1307, ZN => n1820);
   U1637 : AOI211_X1 port map( C1 => registers_15_22_port, C2 => n4931, A => 
                           n1324, B => n1325, ZN => n1306);
   U1638 : AOI221_X1 port map( B1 => registers_29_22_port, B2 => n4898, C1 => 
                           registers_10_22_port, C2 => n4895, A => n1334, ZN =>
                           n1304);
   U1639 : AOI221_X1 port map( B1 => registers_27_22_port, B2 => n4910, C1 => 
                           registers_7_22_port, C2 => n4907, A => n1331, ZN => 
                           n1305);
   U1640 : NAND4_X1 port map( A1 => n1271, A2 => n1272, A3 => n1273, A4 => 
                           n1274, ZN => n1821);
   U1641 : AOI211_X1 port map( C1 => registers_15_21_port, C2 => n4931, A => 
                           n1291, B => n1292, ZN => n1273);
   U1642 : AOI221_X1 port map( B1 => registers_29_21_port, B2 => n4898, C1 => 
                           registers_10_21_port, C2 => n4895, A => n1301, ZN =>
                           n1271);
   U1643 : AOI221_X1 port map( B1 => registers_27_21_port, B2 => n4910, C1 => 
                           registers_7_21_port, C2 => n4907, A => n1298, ZN => 
                           n1272);
   U1644 : NAND4_X1 port map( A1 => n1238, A2 => n1239, A3 => n1240, A4 => 
                           n1241, ZN => n1822);
   U1645 : AOI211_X1 port map( C1 => registers_15_20_port, C2 => n4931, A => 
                           n1258, B => n1259, ZN => n1240);
   U1646 : AOI221_X1 port map( B1 => registers_29_20_port, B2 => n4898, C1 => 
                           registers_10_20_port, C2 => n4895, A => n1268, ZN =>
                           n1238);
   U1647 : AOI221_X1 port map( B1 => registers_27_20_port, B2 => n4910, C1 => 
                           registers_7_20_port, C2 => n4907, A => n1265, ZN => 
                           n1239);
   U1648 : NAND4_X1 port map( A1 => n1205, A2 => n1206, A3 => n1207, A4 => 
                           n1208, ZN => n1823);
   U1649 : AOI211_X1 port map( C1 => registers_15_19_port, C2 => n4932, A => 
                           n1225, B => n1226, ZN => n1207);
   U1650 : AOI221_X1 port map( B1 => registers_29_19_port, B2 => n4899, C1 => 
                           registers_10_19_port, C2 => n4896, A => n1235, ZN =>
                           n1205);
   U1651 : AOI221_X1 port map( B1 => registers_27_19_port, B2 => n4911, C1 => 
                           registers_7_19_port, C2 => n4908, A => n1232, ZN => 
                           n1206);
   U1652 : NAND4_X1 port map( A1 => n1172, A2 => n1173, A3 => n1174, A4 => 
                           n1175, ZN => n1824);
   U1653 : AOI211_X1 port map( C1 => registers_15_18_port, C2 => n4932, A => 
                           n1192, B => n1193, ZN => n1174);
   U1654 : AOI221_X1 port map( B1 => registers_29_18_port, B2 => n4899, C1 => 
                           registers_10_18_port, C2 => n4896, A => n1202, ZN =>
                           n1172);
   U1655 : AOI221_X1 port map( B1 => registers_27_18_port, B2 => n4911, C1 => 
                           registers_7_18_port, C2 => n4908, A => n1199, ZN => 
                           n1173);
   U1656 : NAND4_X1 port map( A1 => n1139, A2 => n1140, A3 => n1141, A4 => 
                           n1142, ZN => n1825);
   U1657 : AOI211_X1 port map( C1 => registers_15_17_port, C2 => n4932, A => 
                           n1159, B => n1160, ZN => n1141);
   U1658 : AOI221_X1 port map( B1 => registers_29_17_port, B2 => n4899, C1 => 
                           registers_10_17_port, C2 => n4896, A => n1169, ZN =>
                           n1139);
   U1659 : AOI221_X1 port map( B1 => registers_27_17_port, B2 => n4911, C1 => 
                           registers_7_17_port, C2 => n4908, A => n1166, ZN => 
                           n1140);
   U1660 : NAND4_X1 port map( A1 => n1106, A2 => n1107, A3 => n1108, A4 => 
                           n1109, ZN => n1826);
   U1661 : AOI211_X1 port map( C1 => registers_15_16_port, C2 => n4932, A => 
                           n1126, B => n1127, ZN => n1108);
   U1662 : AOI221_X1 port map( B1 => registers_29_16_port, B2 => n4899, C1 => 
                           registers_10_16_port, C2 => n4896, A => n1136, ZN =>
                           n1106);
   U1663 : AOI221_X1 port map( B1 => registers_27_16_port, B2 => n4911, C1 => 
                           registers_7_16_port, C2 => n4908, A => n1133, ZN => 
                           n1107);
   U1664 : NAND2_X1 port map( A1 => r_signal_port_b, A2 => enable, ZN => n3072)
                           ;
   U1665 : NAND2_X1 port map( A1 => r_signal_port_a, A2 => enable, ZN => n3075)
                           ;
   U1666 : INV_X1 port map( A => address_port_b(2), ZN => n2306);
   U1667 : INV_X1 port map( A => address_port_b(1), ZN => n2305);
   U1668 : INV_X1 port map( A => address_port_a(1), ZN => n1649);
   U1669 : INV_X1 port map( A => address_port_a(2), ZN => n1650);
   U1670 : INV_X1 port map( A => address_port_w(2), ZN => n545);
   U1671 : INV_X1 port map( A => address_port_w(0), ZN => n546);
   U1672 : INV_X1 port map( A => address_port_w(1), ZN => n544);
   U1673 : INV_X1 port map( A => registers_31_15_port, ZN => n1081);
   U1674 : INV_X1 port map( A => registers_5_15_port, ZN => n1084);
   U1675 : INV_X1 port map( A => registers_4_15_port, ZN => n1087);
   U1676 : INV_X1 port map( A => registers_16_15_port, ZN => n1090);
   U1677 : INV_X1 port map( A => registers_11_15_port, ZN => n1097);
   U1678 : INV_X1 port map( A => registers_31_14_port, ZN => n1048);
   U1679 : INV_X1 port map( A => registers_5_14_port, ZN => n1051);
   U1680 : INV_X1 port map( A => registers_4_14_port, ZN => n1054);
   U1681 : INV_X1 port map( A => registers_16_14_port, ZN => n1057);
   U1682 : INV_X1 port map( A => registers_11_14_port, ZN => n1064);
   U1683 : INV_X1 port map( A => registers_31_13_port, ZN => n1015);
   U1684 : INV_X1 port map( A => registers_5_13_port, ZN => n1018);
   U1685 : INV_X1 port map( A => registers_4_13_port, ZN => n1021);
   U1686 : INV_X1 port map( A => registers_16_13_port, ZN => n1024);
   U1687 : INV_X1 port map( A => registers_11_13_port, ZN => n1031);
   U1688 : INV_X1 port map( A => registers_31_12_port, ZN => n982);
   U1689 : INV_X1 port map( A => registers_5_12_port, ZN => n985);
   U1690 : INV_X1 port map( A => registers_4_12_port, ZN => n988);
   U1691 : INV_X1 port map( A => registers_16_12_port, ZN => n991);
   U1692 : INV_X1 port map( A => registers_11_12_port, ZN => n998);
   U1693 : INV_X1 port map( A => registers_31_11_port, ZN => n949);
   U1694 : INV_X1 port map( A => registers_5_11_port, ZN => n952);
   U1695 : INV_X1 port map( A => registers_4_11_port, ZN => n955);
   U1696 : INV_X1 port map( A => registers_16_11_port, ZN => n958);
   U1697 : INV_X1 port map( A => registers_11_11_port, ZN => n965);
   U1698 : INV_X1 port map( A => registers_31_10_port, ZN => n916);
   U1699 : INV_X1 port map( A => registers_5_10_port, ZN => n919);
   U1700 : INV_X1 port map( A => registers_4_10_port, ZN => n922);
   U1701 : INV_X1 port map( A => registers_16_10_port, ZN => n925);
   U1702 : INV_X1 port map( A => registers_11_10_port, ZN => n932);
   U1703 : INV_X1 port map( A => registers_31_9_port, ZN => n883);
   U1704 : INV_X1 port map( A => registers_5_9_port, ZN => n886);
   U1705 : INV_X1 port map( A => registers_4_9_port, ZN => n889);
   U1706 : INV_X1 port map( A => registers_16_9_port, ZN => n892);
   U1707 : INV_X1 port map( A => registers_11_9_port, ZN => n899);
   U1708 : INV_X1 port map( A => registers_31_8_port, ZN => n850);
   U1709 : INV_X1 port map( A => registers_5_8_port, ZN => n853);
   U1710 : INV_X1 port map( A => registers_4_8_port, ZN => n856);
   U1711 : INV_X1 port map( A => registers_16_8_port, ZN => n859);
   U1712 : INV_X1 port map( A => registers_11_8_port, ZN => n866);
   U1713 : INV_X1 port map( A => registers_31_7_port, ZN => n817);
   U1714 : INV_X1 port map( A => registers_5_7_port, ZN => n820);
   U1715 : INV_X1 port map( A => registers_4_7_port, ZN => n823);
   U1716 : INV_X1 port map( A => registers_16_7_port, ZN => n826);
   U1717 : INV_X1 port map( A => registers_11_7_port, ZN => n833);
   U1718 : INV_X1 port map( A => registers_31_6_port, ZN => n784);
   U1719 : INV_X1 port map( A => registers_5_6_port, ZN => n787);
   U1720 : INV_X1 port map( A => registers_4_6_port, ZN => n790);
   U1721 : INV_X1 port map( A => registers_16_6_port, ZN => n793);
   U1722 : INV_X1 port map( A => registers_11_6_port, ZN => n800);
   U1723 : INV_X1 port map( A => registers_31_5_port, ZN => n751);
   U1724 : INV_X1 port map( A => registers_5_5_port, ZN => n754);
   U1725 : INV_X1 port map( A => registers_4_5_port, ZN => n757);
   U1726 : INV_X1 port map( A => registers_16_5_port, ZN => n760);
   U1727 : INV_X1 port map( A => registers_11_5_port, ZN => n767);
   U1728 : INV_X1 port map( A => registers_31_4_port, ZN => n718);
   U1729 : INV_X1 port map( A => registers_5_4_port, ZN => n721);
   U1730 : INV_X1 port map( A => registers_4_4_port, ZN => n724);
   U1731 : INV_X1 port map( A => registers_16_4_port, ZN => n727);
   U1732 : INV_X1 port map( A => registers_11_4_port, ZN => n734);
   U1733 : INV_X1 port map( A => registers_31_3_port, ZN => n685);
   U1734 : INV_X1 port map( A => registers_5_3_port, ZN => n688);
   U1735 : INV_X1 port map( A => registers_4_3_port, ZN => n691);
   U1736 : INV_X1 port map( A => registers_16_3_port, ZN => n694);
   U1737 : INV_X1 port map( A => registers_11_3_port, ZN => n701);
   U1738 : INV_X1 port map( A => registers_31_2_port, ZN => n652);
   U1739 : INV_X1 port map( A => registers_5_2_port, ZN => n655);
   U1740 : INV_X1 port map( A => registers_4_2_port, ZN => n658);
   U1741 : INV_X1 port map( A => registers_16_2_port, ZN => n661);
   U1742 : INV_X1 port map( A => registers_11_2_port, ZN => n668);
   U1743 : INV_X1 port map( A => registers_31_1_port, ZN => n619);
   U1744 : INV_X1 port map( A => registers_5_1_port, ZN => n622);
   U1745 : INV_X1 port map( A => registers_4_1_port, ZN => n625);
   U1746 : INV_X1 port map( A => registers_16_1_port, ZN => n628);
   U1747 : INV_X1 port map( A => registers_11_1_port, ZN => n635);
   U1748 : INV_X1 port map( A => registers_31_0_port, ZN => n556);
   U1749 : INV_X1 port map( A => registers_5_0_port, ZN => n563);
   U1750 : INV_X1 port map( A => registers_4_0_port, ZN => n570);
   U1751 : INV_X1 port map( A => registers_16_0_port, ZN => n577);
   U1752 : INV_X1 port map( A => registers_11_0_port, ZN => n591);
   U1753 : INV_X1 port map( A => registers_31_31_port, ZN => n1609);
   U1754 : INV_X1 port map( A => registers_5_31_port, ZN => n1619);
   U1755 : INV_X1 port map( A => registers_4_31_port, ZN => n1625);
   U1756 : INV_X1 port map( A => registers_16_31_port, ZN => n1630);
   U1757 : INV_X1 port map( A => registers_11_31_port, ZN => n1638);
   U1758 : INV_X1 port map( A => registers_31_30_port, ZN => n1576);
   U1759 : INV_X1 port map( A => registers_5_30_port, ZN => n1579);
   U1760 : INV_X1 port map( A => registers_4_30_port, ZN => n1582);
   U1761 : INV_X1 port map( A => registers_16_30_port, ZN => n1585);
   U1762 : INV_X1 port map( A => registers_11_30_port, ZN => n1592);
   U1763 : INV_X1 port map( A => registers_31_29_port, ZN => n1543);
   U1764 : INV_X1 port map( A => registers_5_29_port, ZN => n1546);
   U1765 : INV_X1 port map( A => registers_4_29_port, ZN => n1549);
   U1766 : INV_X1 port map( A => registers_16_29_port, ZN => n1552);
   U1767 : INV_X1 port map( A => registers_11_29_port, ZN => n1559);
   U1768 : INV_X1 port map( A => registers_31_28_port, ZN => n1510);
   U1769 : INV_X1 port map( A => registers_5_28_port, ZN => n1513);
   U1770 : INV_X1 port map( A => registers_4_28_port, ZN => n1516);
   U1771 : INV_X1 port map( A => registers_16_28_port, ZN => n1519);
   U1772 : INV_X1 port map( A => registers_11_28_port, ZN => n1526);
   U1773 : INV_X1 port map( A => registers_31_27_port, ZN => n1477);
   U1774 : INV_X1 port map( A => registers_5_27_port, ZN => n1480);
   U1775 : INV_X1 port map( A => registers_4_27_port, ZN => n1483);
   U1776 : INV_X1 port map( A => registers_16_27_port, ZN => n1486);
   U1777 : INV_X1 port map( A => registers_11_27_port, ZN => n1493);
   U1778 : INV_X1 port map( A => registers_31_26_port, ZN => n1444);
   U1779 : INV_X1 port map( A => registers_5_26_port, ZN => n1447);
   U1780 : INV_X1 port map( A => registers_4_26_port, ZN => n1450);
   U1781 : INV_X1 port map( A => registers_16_26_port, ZN => n1453);
   U1782 : INV_X1 port map( A => registers_11_26_port, ZN => n1460);
   U1783 : INV_X1 port map( A => registers_31_25_port, ZN => n1411);
   U1784 : INV_X1 port map( A => registers_5_25_port, ZN => n1414);
   U1785 : INV_X1 port map( A => registers_4_25_port, ZN => n1417);
   U1786 : INV_X1 port map( A => registers_16_25_port, ZN => n1420);
   U1787 : INV_X1 port map( A => registers_11_25_port, ZN => n1427);
   U1788 : INV_X1 port map( A => registers_31_24_port, ZN => n1378);
   U1789 : INV_X1 port map( A => registers_5_24_port, ZN => n1381);
   U1790 : INV_X1 port map( A => registers_4_24_port, ZN => n1384);
   U1791 : INV_X1 port map( A => registers_16_24_port, ZN => n1387);
   U1792 : INV_X1 port map( A => registers_11_24_port, ZN => n1394);
   U1793 : INV_X1 port map( A => registers_31_23_port, ZN => n1345);
   U1794 : INV_X1 port map( A => registers_5_23_port, ZN => n1348);
   U1795 : INV_X1 port map( A => registers_4_23_port, ZN => n1351);
   U1796 : INV_X1 port map( A => registers_16_23_port, ZN => n1354);
   U1797 : INV_X1 port map( A => registers_11_23_port, ZN => n1361);
   U1798 : INV_X1 port map( A => registers_31_22_port, ZN => n1312);
   U1799 : INV_X1 port map( A => registers_5_22_port, ZN => n1315);
   U1800 : INV_X1 port map( A => registers_4_22_port, ZN => n1318);
   U1801 : INV_X1 port map( A => registers_16_22_port, ZN => n1321);
   U1802 : INV_X1 port map( A => registers_11_22_port, ZN => n1328);
   U1803 : INV_X1 port map( A => registers_31_21_port, ZN => n1279);
   U1804 : INV_X1 port map( A => registers_5_21_port, ZN => n1282);
   U1805 : INV_X1 port map( A => registers_4_21_port, ZN => n1285);
   U1806 : INV_X1 port map( A => registers_16_21_port, ZN => n1288);
   U1807 : INV_X1 port map( A => registers_11_21_port, ZN => n1295);
   U1808 : INV_X1 port map( A => registers_31_20_port, ZN => n1246);
   U1809 : INV_X1 port map( A => registers_5_20_port, ZN => n1249);
   U1810 : INV_X1 port map( A => registers_4_20_port, ZN => n1252);
   U1811 : INV_X1 port map( A => registers_16_20_port, ZN => n1255);
   U1812 : INV_X1 port map( A => registers_11_20_port, ZN => n1262);
   U1813 : INV_X1 port map( A => registers_31_19_port, ZN => n1213);
   U1814 : INV_X1 port map( A => registers_5_19_port, ZN => n1216);
   U1815 : INV_X1 port map( A => registers_4_19_port, ZN => n1219);
   U1816 : INV_X1 port map( A => registers_16_19_port, ZN => n1222);
   U1817 : INV_X1 port map( A => registers_11_19_port, ZN => n1229);
   U1818 : INV_X1 port map( A => registers_31_18_port, ZN => n1180);
   U1819 : INV_X1 port map( A => registers_5_18_port, ZN => n1183);
   U1820 : INV_X1 port map( A => registers_4_18_port, ZN => n1186);
   U1821 : INV_X1 port map( A => registers_16_18_port, ZN => n1189);
   U1822 : INV_X1 port map( A => registers_11_18_port, ZN => n1196);
   U1823 : INV_X1 port map( A => registers_31_17_port, ZN => n1147);
   U1824 : INV_X1 port map( A => registers_5_17_port, ZN => n1150);
   U1825 : INV_X1 port map( A => registers_4_17_port, ZN => n1153);
   U1826 : INV_X1 port map( A => registers_16_17_port, ZN => n1156);
   U1827 : INV_X1 port map( A => registers_11_17_port, ZN => n1163);
   U1828 : INV_X1 port map( A => registers_31_16_port, ZN => n1114);
   U1829 : INV_X1 port map( A => registers_5_16_port, ZN => n1117);
   U1830 : INV_X1 port map( A => registers_4_16_port, ZN => n1120);
   U1831 : INV_X1 port map( A => registers_16_16_port, ZN => n1123);
   U1832 : INV_X1 port map( A => registers_11_16_port, ZN => n1130);
   U1833 : INV_X1 port map( A => registers_6_15_port, ZN => n1101);
   U1846 : INV_X1 port map( A => registers_23_15_port, ZN => n1104);
   U1847 : INV_X1 port map( A => registers_22_15_port, ZN => n1095);
   U1848 : INV_X1 port map( A => registers_6_14_port, ZN => n1068);
   U1849 : INV_X1 port map( A => registers_23_14_port, ZN => n1071);
   U1850 : INV_X1 port map( A => registers_22_14_port, ZN => n1062);
   U1851 : INV_X1 port map( A => registers_6_13_port, ZN => n1035);
   U1852 : INV_X1 port map( A => registers_23_13_port, ZN => n1038);
   U1853 : INV_X1 port map( A => registers_22_13_port, ZN => n1029);
   U1854 : INV_X1 port map( A => registers_6_12_port, ZN => n1002);
   U1855 : INV_X1 port map( A => registers_23_12_port, ZN => n1005);
   U1856 : INV_X1 port map( A => registers_22_12_port, ZN => n996);
   U1857 : INV_X1 port map( A => registers_6_11_port, ZN => n969);
   U1858 : INV_X1 port map( A => registers_23_11_port, ZN => n972);
   U1859 : INV_X1 port map( A => registers_22_11_port, ZN => n963);
   U1860 : INV_X1 port map( A => registers_6_10_port, ZN => n936);
   U1861 : INV_X1 port map( A => registers_23_10_port, ZN => n939);
   U1862 : INV_X1 port map( A => registers_22_10_port, ZN => n930);
   U1863 : INV_X1 port map( A => registers_6_9_port, ZN => n903);
   U1864 : INV_X1 port map( A => registers_23_9_port, ZN => n906);
   U1865 : INV_X1 port map( A => registers_22_9_port, ZN => n897);
   U1866 : INV_X1 port map( A => registers_6_8_port, ZN => n870);
   U1867 : INV_X1 port map( A => registers_23_8_port, ZN => n873);
   U1868 : INV_X1 port map( A => registers_22_8_port, ZN => n864);
   U1869 : INV_X1 port map( A => registers_6_7_port, ZN => n837);
   U1870 : INV_X1 port map( A => registers_23_7_port, ZN => n840);
   U1871 : INV_X1 port map( A => registers_22_7_port, ZN => n831);
   U1872 : INV_X1 port map( A => registers_6_6_port, ZN => n804);
   U1873 : INV_X1 port map( A => registers_23_6_port, ZN => n807);
   U1874 : INV_X1 port map( A => registers_22_6_port, ZN => n798);
   U1875 : INV_X1 port map( A => registers_6_5_port, ZN => n771);
   U1876 : INV_X1 port map( A => registers_23_5_port, ZN => n774);
   U1877 : INV_X1 port map( A => registers_22_5_port, ZN => n765);
   U1878 : INV_X1 port map( A => registers_6_4_port, ZN => n738);
   U1879 : INV_X1 port map( A => registers_23_4_port, ZN => n741);
   U1880 : INV_X1 port map( A => registers_22_4_port, ZN => n732);
   U1881 : INV_X1 port map( A => registers_6_3_port, ZN => n705);
   U1882 : INV_X1 port map( A => registers_23_3_port, ZN => n708);
   U1883 : INV_X1 port map( A => registers_22_3_port, ZN => n699);
   U1884 : INV_X1 port map( A => registers_6_2_port, ZN => n672);
   U1885 : INV_X1 port map( A => registers_23_2_port, ZN => n675);
   U1886 : INV_X1 port map( A => registers_22_2_port, ZN => n666);
   U1887 : INV_X1 port map( A => registers_6_1_port, ZN => n639);
   U1888 : INV_X1 port map( A => registers_23_1_port, ZN => n642);
   U1889 : INV_X1 port map( A => registers_22_1_port, ZN => n633);
   U1890 : INV_X1 port map( A => registers_6_0_port, ZN => n601);
   U1891 : INV_X1 port map( A => registers_23_0_port, ZN => n608);
   U1892 : INV_X1 port map( A => registers_22_0_port, ZN => n587);
   U1893 : INV_X1 port map( A => registers_6_31_port, ZN => n1644);
   U1894 : INV_X1 port map( A => registers_23_31_port, ZN => n1647);
   U1895 : INV_X1 port map( A => registers_22_31_port, ZN => n1635);
   U1896 : INV_X1 port map( A => registers_6_30_port, ZN => n1596);
   U1897 : INV_X1 port map( A => registers_23_30_port, ZN => n1599);
   U1898 : INV_X1 port map( A => registers_22_30_port, ZN => n1590);
   U1899 : INV_X1 port map( A => registers_6_29_port, ZN => n1563);
   U1900 : INV_X1 port map( A => registers_23_29_port, ZN => n1566);
   U1901 : INV_X1 port map( A => registers_22_29_port, ZN => n1557);
   U1902 : INV_X1 port map( A => registers_6_28_port, ZN => n1530);
   U1903 : INV_X1 port map( A => registers_23_28_port, ZN => n1533);
   U1904 : INV_X1 port map( A => registers_22_28_port, ZN => n1524);
   U1905 : INV_X1 port map( A => registers_6_27_port, ZN => n1497);
   U1906 : INV_X1 port map( A => registers_23_27_port, ZN => n1500);
   U1907 : INV_X1 port map( A => registers_22_27_port, ZN => n1491);
   U1908 : INV_X1 port map( A => registers_6_26_port, ZN => n1464);
   U1909 : INV_X1 port map( A => registers_23_26_port, ZN => n1467);
   U1910 : INV_X1 port map( A => registers_22_26_port, ZN => n1458);
   U1911 : INV_X1 port map( A => registers_6_25_port, ZN => n1431);
   U1912 : INV_X1 port map( A => registers_23_25_port, ZN => n1434);
   U1913 : INV_X1 port map( A => registers_22_25_port, ZN => n1425);
   U1914 : INV_X1 port map( A => registers_6_24_port, ZN => n1398);
   U1915 : INV_X1 port map( A => registers_23_24_port, ZN => n1401);
   U1916 : INV_X1 port map( A => registers_22_24_port, ZN => n1392);
   U1917 : INV_X1 port map( A => registers_6_23_port, ZN => n1365);
   U1918 : INV_X1 port map( A => registers_23_23_port, ZN => n1368);
   U1919 : INV_X1 port map( A => registers_22_23_port, ZN => n1359);
   U1920 : INV_X1 port map( A => registers_6_22_port, ZN => n1332);
   U1921 : INV_X1 port map( A => registers_23_22_port, ZN => n1335);
   U1922 : INV_X1 port map( A => registers_22_22_port, ZN => n1326);
   U1923 : INV_X1 port map( A => registers_6_21_port, ZN => n1299);
   U1924 : INV_X1 port map( A => registers_23_21_port, ZN => n1302);
   U1925 : INV_X1 port map( A => registers_22_21_port, ZN => n1293);
   U1926 : INV_X1 port map( A => registers_6_20_port, ZN => n1266);
   U1927 : INV_X1 port map( A => registers_23_20_port, ZN => n1269);
   U1928 : INV_X1 port map( A => registers_22_20_port, ZN => n1260);
   U1929 : INV_X1 port map( A => registers_6_19_port, ZN => n1233);
   U1930 : INV_X1 port map( A => registers_23_19_port, ZN => n1236);
   U1931 : INV_X1 port map( A => registers_22_19_port, ZN => n1227);
   U1932 : INV_X1 port map( A => registers_6_18_port, ZN => n1200);
   U1933 : INV_X1 port map( A => registers_23_18_port, ZN => n1203);
   U1934 : INV_X1 port map( A => registers_22_18_port, ZN => n1194);
   U1935 : INV_X1 port map( A => registers_6_17_port, ZN => n1167);
   U1936 : INV_X1 port map( A => registers_23_17_port, ZN => n1170);
   U1937 : INV_X1 port map( A => registers_22_17_port, ZN => n1161);
   U1938 : INV_X1 port map( A => registers_6_16_port, ZN => n1134);
   U1939 : INV_X1 port map( A => registers_23_16_port, ZN => n1137);
   U1940 : INV_X1 port map( A => registers_22_16_port, ZN => n1128);
   U1941 : INV_X1 port map( A => registers_2_15_port, ZN => n1102);
   U1942 : INV_X1 port map( A => registers_26_15_port, ZN => n1105);
   U1943 : INV_X1 port map( A => registers_19_15_port, ZN => n1096);
   U1944 : INV_X1 port map( A => registers_2_14_port, ZN => n1069);
   U1945 : INV_X1 port map( A => registers_26_14_port, ZN => n1072);
   U1946 : INV_X1 port map( A => registers_19_14_port, ZN => n1063);
   U1947 : INV_X1 port map( A => registers_2_13_port, ZN => n1036);
   U1948 : INV_X1 port map( A => registers_26_13_port, ZN => n1039);
   U1949 : INV_X1 port map( A => registers_19_13_port, ZN => n1030);
   U1950 : INV_X1 port map( A => registers_2_12_port, ZN => n1003);
   U1951 : INV_X1 port map( A => registers_26_12_port, ZN => n1006);
   U1952 : INV_X1 port map( A => registers_19_12_port, ZN => n997);
   U1953 : INV_X1 port map( A => registers_2_11_port, ZN => n970);
   U1954 : INV_X1 port map( A => registers_26_11_port, ZN => n973);
   U1955 : INV_X1 port map( A => registers_19_11_port, ZN => n964);
   U1956 : INV_X1 port map( A => registers_2_10_port, ZN => n937);
   U1957 : INV_X1 port map( A => registers_26_10_port, ZN => n940);
   U1958 : INV_X1 port map( A => registers_19_10_port, ZN => n931);
   U1959 : INV_X1 port map( A => registers_2_9_port, ZN => n904);
   U1960 : INV_X1 port map( A => registers_26_9_port, ZN => n907);
   U1961 : INV_X1 port map( A => registers_19_9_port, ZN => n898);
   U1962 : INV_X1 port map( A => registers_2_8_port, ZN => n871);
   U1963 : INV_X1 port map( A => registers_26_8_port, ZN => n874);
   U1964 : INV_X1 port map( A => registers_19_8_port, ZN => n865);
   U1965 : INV_X1 port map( A => registers_2_7_port, ZN => n838);
   U1966 : INV_X1 port map( A => registers_26_7_port, ZN => n841);
   U1967 : INV_X1 port map( A => registers_19_7_port, ZN => n832);
   U1968 : INV_X1 port map( A => registers_2_6_port, ZN => n805);
   U1969 : INV_X1 port map( A => registers_26_6_port, ZN => n808);
   U1970 : INV_X1 port map( A => registers_19_6_port, ZN => n799);
   U1971 : INV_X1 port map( A => registers_2_5_port, ZN => n772);
   U1972 : INV_X1 port map( A => registers_26_5_port, ZN => n775);
   U1973 : INV_X1 port map( A => registers_19_5_port, ZN => n766);
   U1974 : INV_X1 port map( A => registers_2_4_port, ZN => n739);
   U1975 : INV_X1 port map( A => registers_26_4_port, ZN => n742);
   U1976 : INV_X1 port map( A => registers_19_4_port, ZN => n733);
   U1977 : INV_X1 port map( A => registers_2_3_port, ZN => n706);
   U1978 : INV_X1 port map( A => registers_26_3_port, ZN => n709);
   U1979 : INV_X1 port map( A => registers_19_3_port, ZN => n700);
   U1980 : INV_X1 port map( A => registers_2_2_port, ZN => n673);
   U1981 : INV_X1 port map( A => registers_26_2_port, ZN => n676);
   U1982 : INV_X1 port map( A => registers_19_2_port, ZN => n667);
   U1983 : INV_X1 port map( A => registers_2_1_port, ZN => n640);
   U1984 : INV_X1 port map( A => registers_26_1_port, ZN => n643);
   U1985 : INV_X1 port map( A => registers_19_1_port, ZN => n634);
   U1986 : INV_X1 port map( A => registers_2_0_port, ZN => n603);
   U1987 : INV_X1 port map( A => registers_26_0_port, ZN => n610);
   U1988 : INV_X1 port map( A => registers_19_0_port, ZN => n589);
   U1989 : INV_X1 port map( A => registers_2_31_port, ZN => n1645);
   U1990 : INV_X1 port map( A => registers_26_31_port, ZN => n1648);
   U1991 : INV_X1 port map( A => registers_19_31_port, ZN => n1636);
   U1992 : INV_X1 port map( A => registers_2_30_port, ZN => n1597);
   U1993 : INV_X1 port map( A => registers_26_30_port, ZN => n1600);
   U1994 : INV_X1 port map( A => registers_19_30_port, ZN => n1591);
   U1995 : INV_X1 port map( A => registers_2_29_port, ZN => n1564);
   U1996 : INV_X1 port map( A => registers_26_29_port, ZN => n1567);
   U1997 : INV_X1 port map( A => registers_19_29_port, ZN => n1558);
   U1998 : INV_X1 port map( A => registers_2_28_port, ZN => n1531);
   U1999 : INV_X1 port map( A => registers_26_28_port, ZN => n1534);
   U2000 : INV_X1 port map( A => registers_19_28_port, ZN => n1525);
   U2001 : INV_X1 port map( A => registers_2_27_port, ZN => n1498);
   U2002 : INV_X1 port map( A => registers_26_27_port, ZN => n1501);
   U2003 : INV_X1 port map( A => registers_19_27_port, ZN => n1492);
   U2004 : INV_X1 port map( A => registers_2_26_port, ZN => n1465);
   U2005 : INV_X1 port map( A => registers_26_26_port, ZN => n1468);
   U2006 : INV_X1 port map( A => registers_19_26_port, ZN => n1459);
   U2007 : INV_X1 port map( A => registers_2_25_port, ZN => n1432);
   U2008 : INV_X1 port map( A => registers_26_25_port, ZN => n1435);
   U2009 : INV_X1 port map( A => registers_19_25_port, ZN => n1426);
   U2010 : INV_X1 port map( A => registers_2_24_port, ZN => n1399);
   U2011 : INV_X1 port map( A => registers_26_24_port, ZN => n1402);
   U2012 : INV_X1 port map( A => registers_19_24_port, ZN => n1393);
   U2013 : INV_X1 port map( A => registers_2_23_port, ZN => n1366);
   U2014 : INV_X1 port map( A => registers_26_23_port, ZN => n1369);
   U2015 : INV_X1 port map( A => registers_19_23_port, ZN => n1360);
   U2016 : INV_X1 port map( A => registers_2_22_port, ZN => n1333);
   U2017 : INV_X1 port map( A => registers_26_22_port, ZN => n1336);
   U2018 : INV_X1 port map( A => registers_19_22_port, ZN => n1327);
   U2019 : INV_X1 port map( A => registers_2_21_port, ZN => n1300);
   U2020 : INV_X1 port map( A => registers_26_21_port, ZN => n1303);
   U2021 : INV_X1 port map( A => registers_19_21_port, ZN => n1294);
   U2022 : INV_X1 port map( A => registers_2_20_port, ZN => n1267);
   U2023 : INV_X1 port map( A => registers_26_20_port, ZN => n1270);
   U2024 : INV_X1 port map( A => registers_19_20_port, ZN => n1261);
   U2025 : INV_X1 port map( A => registers_2_19_port, ZN => n1234);
   U2026 : INV_X1 port map( A => registers_26_19_port, ZN => n1237);
   U2027 : INV_X1 port map( A => registers_19_19_port, ZN => n1228);
   U2028 : INV_X1 port map( A => registers_2_18_port, ZN => n1201);
   U2029 : INV_X1 port map( A => registers_26_18_port, ZN => n1204);
   U2030 : INV_X1 port map( A => registers_19_18_port, ZN => n1195);
   U2031 : INV_X1 port map( A => registers_2_17_port, ZN => n1168);
   U2032 : INV_X1 port map( A => registers_26_17_port, ZN => n1171);
   U2033 : INV_X1 port map( A => registers_19_17_port, ZN => n1162);
   U2034 : INV_X1 port map( A => registers_2_16_port, ZN => n1135);
   U2035 : INV_X1 port map( A => registers_26_16_port, ZN => n1138);
   U2036 : INV_X1 port map( A => registers_19_16_port, ZN => n1129);
   U2037 : INV_X1 port map( A => registers_9_15_port, ZN => n1082);
   U2038 : INV_X1 port map( A => registers_8_15_port, ZN => n1085);
   U2039 : INV_X1 port map( A => registers_1_15_port, ZN => n1088);
   U2040 : INV_X1 port map( A => registers_17_15_port, ZN => n1091);
   U2041 : INV_X1 port map( A => registers_3_15_port, ZN => n1098);
   U2042 : INV_X1 port map( A => registers_9_14_port, ZN => n1049);
   U2043 : INV_X1 port map( A => registers_8_14_port, ZN => n1052);
   U2044 : INV_X1 port map( A => registers_1_14_port, ZN => n1055);
   U2045 : INV_X1 port map( A => registers_17_14_port, ZN => n1058);
   U2046 : INV_X1 port map( A => registers_3_14_port, ZN => n1065);
   U2047 : INV_X1 port map( A => registers_9_13_port, ZN => n1016);
   U2048 : INV_X1 port map( A => registers_8_13_port, ZN => n1019);
   U2049 : INV_X1 port map( A => registers_1_13_port, ZN => n1022);
   U2050 : INV_X1 port map( A => registers_17_13_port, ZN => n1025);
   U2051 : INV_X1 port map( A => registers_3_13_port, ZN => n1032);
   U2052 : INV_X1 port map( A => registers_9_12_port, ZN => n983);
   U2053 : INV_X1 port map( A => registers_8_12_port, ZN => n986);
   U2054 : INV_X1 port map( A => registers_1_12_port, ZN => n989);
   U2055 : INV_X1 port map( A => registers_17_12_port, ZN => n992);
   U2056 : INV_X1 port map( A => registers_3_12_port, ZN => n999);
   U2057 : INV_X1 port map( A => registers_9_11_port, ZN => n950);
   U2058 : INV_X1 port map( A => registers_8_11_port, ZN => n953);
   U2059 : INV_X1 port map( A => registers_1_11_port, ZN => n956);
   U2060 : INV_X1 port map( A => registers_17_11_port, ZN => n959);
   U2061 : INV_X1 port map( A => registers_3_11_port, ZN => n966);
   U2062 : INV_X1 port map( A => registers_9_10_port, ZN => n917);
   U2063 : INV_X1 port map( A => registers_8_10_port, ZN => n920);
   U2064 : INV_X1 port map( A => registers_1_10_port, ZN => n923);
   U2065 : INV_X1 port map( A => registers_17_10_port, ZN => n926);
   U2066 : INV_X1 port map( A => registers_3_10_port, ZN => n933);
   U2067 : INV_X1 port map( A => registers_9_9_port, ZN => n884);
   U2068 : INV_X1 port map( A => registers_8_9_port, ZN => n887);
   U2069 : INV_X1 port map( A => registers_1_9_port, ZN => n890);
   U2070 : INV_X1 port map( A => registers_17_9_port, ZN => n893);
   U2071 : INV_X1 port map( A => registers_3_9_port, ZN => n900);
   U2072 : INV_X1 port map( A => registers_9_8_port, ZN => n851);
   U2073 : INV_X1 port map( A => registers_8_8_port, ZN => n854);
   U2074 : INV_X1 port map( A => registers_1_8_port, ZN => n857);
   U2075 : INV_X1 port map( A => registers_17_8_port, ZN => n860);
   U2076 : INV_X1 port map( A => registers_3_8_port, ZN => n867);
   U2077 : INV_X1 port map( A => registers_9_7_port, ZN => n818);
   U2078 : INV_X1 port map( A => registers_8_7_port, ZN => n821);
   U2079 : INV_X1 port map( A => registers_1_7_port, ZN => n824);
   U2080 : INV_X1 port map( A => registers_17_7_port, ZN => n827);
   U2081 : INV_X1 port map( A => registers_3_7_port, ZN => n834);
   U2082 : INV_X1 port map( A => registers_9_6_port, ZN => n785);
   U2083 : INV_X1 port map( A => registers_8_6_port, ZN => n788);
   U2084 : INV_X1 port map( A => registers_1_6_port, ZN => n791);
   U2085 : INV_X1 port map( A => registers_17_6_port, ZN => n794);
   U2086 : INV_X1 port map( A => registers_3_6_port, ZN => n801);
   U2087 : INV_X1 port map( A => registers_9_5_port, ZN => n752);
   U2088 : INV_X1 port map( A => registers_8_5_port, ZN => n755);
   U2089 : INV_X1 port map( A => registers_1_5_port, ZN => n758);
   U2090 : INV_X1 port map( A => registers_17_5_port, ZN => n761);
   U2091 : INV_X1 port map( A => registers_3_5_port, ZN => n768);
   U2092 : INV_X1 port map( A => registers_9_4_port, ZN => n719);
   U2093 : INV_X1 port map( A => registers_8_4_port, ZN => n722);
   U2094 : INV_X1 port map( A => registers_1_4_port, ZN => n725);
   U2095 : INV_X1 port map( A => registers_17_4_port, ZN => n728);
   U2096 : INV_X1 port map( A => registers_3_4_port, ZN => n735);
   U2097 : INV_X1 port map( A => registers_9_3_port, ZN => n686);
   U2098 : INV_X1 port map( A => registers_8_3_port, ZN => n689);
   U2099 : INV_X1 port map( A => registers_1_3_port, ZN => n692);
   U2100 : INV_X1 port map( A => registers_17_3_port, ZN => n695);
   U2101 : INV_X1 port map( A => registers_3_3_port, ZN => n702);
   U2102 : INV_X1 port map( A => registers_9_2_port, ZN => n653);
   U2103 : INV_X1 port map( A => registers_8_2_port, ZN => n656);
   U2104 : INV_X1 port map( A => registers_1_2_port, ZN => n659);
   U2105 : INV_X1 port map( A => registers_17_2_port, ZN => n662);
   U2106 : INV_X1 port map( A => registers_3_2_port, ZN => n669);
   U2107 : INV_X1 port map( A => registers_9_1_port, ZN => n620);
   U2108 : INV_X1 port map( A => registers_8_1_port, ZN => n623);
   U2109 : INV_X1 port map( A => registers_1_1_port, ZN => n626);
   U2110 : INV_X1 port map( A => registers_17_1_port, ZN => n629);
   U2111 : INV_X1 port map( A => registers_3_1_port, ZN => n636);
   U2112 : INV_X1 port map( A => registers_9_0_port, ZN => n558);
   U2113 : INV_X1 port map( A => registers_8_0_port, ZN => n565);
   U2114 : INV_X1 port map( A => registers_1_0_port, ZN => n572);
   U2115 : INV_X1 port map( A => registers_17_0_port, ZN => n579);
   U2116 : INV_X1 port map( A => registers_3_0_port, ZN => n593);
   U2117 : INV_X1 port map( A => registers_9_31_port, ZN => n1610);
   U2118 : INV_X1 port map( A => registers_8_31_port, ZN => n1620);
   U2119 : INV_X1 port map( A => registers_1_31_port, ZN => n1626);
   U2120 : INV_X1 port map( A => registers_17_31_port, ZN => n1631);
   U2121 : INV_X1 port map( A => registers_3_31_port, ZN => n1639);
   U2122 : INV_X1 port map( A => registers_9_30_port, ZN => n1577);
   U2123 : INV_X1 port map( A => registers_8_30_port, ZN => n1580);
   U2124 : INV_X1 port map( A => registers_1_30_port, ZN => n1583);
   U2125 : INV_X1 port map( A => registers_17_30_port, ZN => n1586);
   U2126 : INV_X1 port map( A => registers_3_30_port, ZN => n1593);
   U2127 : INV_X1 port map( A => registers_9_29_port, ZN => n1544);
   U2128 : INV_X1 port map( A => registers_8_29_port, ZN => n1547);
   U2129 : INV_X1 port map( A => registers_1_29_port, ZN => n1550);
   U2130 : INV_X1 port map( A => registers_17_29_port, ZN => n1553);
   U2131 : INV_X1 port map( A => registers_3_29_port, ZN => n1560);
   U2132 : INV_X1 port map( A => registers_9_28_port, ZN => n1511);
   U2133 : INV_X1 port map( A => registers_8_28_port, ZN => n1514);
   U2134 : INV_X1 port map( A => registers_1_28_port, ZN => n1517);
   U2135 : INV_X1 port map( A => registers_17_28_port, ZN => n1520);
   U2136 : INV_X1 port map( A => registers_3_28_port, ZN => n1527);
   U2137 : INV_X1 port map( A => registers_9_27_port, ZN => n1478);
   U2138 : INV_X1 port map( A => registers_8_27_port, ZN => n1481);
   U2139 : INV_X1 port map( A => registers_1_27_port, ZN => n1484);
   U2140 : INV_X1 port map( A => registers_17_27_port, ZN => n1487);
   U2141 : INV_X1 port map( A => registers_3_27_port, ZN => n1494);
   U2142 : INV_X1 port map( A => registers_9_26_port, ZN => n1445);
   U2143 : INV_X1 port map( A => registers_8_26_port, ZN => n1448);
   U2144 : INV_X1 port map( A => registers_1_26_port, ZN => n1451);
   U2145 : INV_X1 port map( A => registers_17_26_port, ZN => n1454);
   U2146 : INV_X1 port map( A => registers_3_26_port, ZN => n1461);
   U2147 : INV_X1 port map( A => registers_9_25_port, ZN => n1412);
   U2148 : INV_X1 port map( A => registers_8_25_port, ZN => n1415);
   U2149 : INV_X1 port map( A => registers_1_25_port, ZN => n1418);
   U2150 : INV_X1 port map( A => registers_17_25_port, ZN => n1421);
   U2151 : INV_X1 port map( A => registers_3_25_port, ZN => n1428);
   U2152 : INV_X1 port map( A => registers_9_24_port, ZN => n1379);
   U2153 : INV_X1 port map( A => registers_8_24_port, ZN => n1382);
   U2154 : INV_X1 port map( A => registers_1_24_port, ZN => n1385);
   U2155 : INV_X1 port map( A => registers_17_24_port, ZN => n1388);
   U2156 : INV_X1 port map( A => registers_3_24_port, ZN => n1395);
   U2157 : INV_X1 port map( A => registers_9_23_port, ZN => n1346);
   U2158 : INV_X1 port map( A => registers_8_23_port, ZN => n1349);
   U2159 : INV_X1 port map( A => registers_1_23_port, ZN => n1352);
   U2160 : INV_X1 port map( A => registers_17_23_port, ZN => n1355);
   U2161 : INV_X1 port map( A => registers_3_23_port, ZN => n1362);
   U2162 : INV_X1 port map( A => registers_9_22_port, ZN => n1313);
   U2163 : INV_X1 port map( A => registers_8_22_port, ZN => n1316);
   U2164 : INV_X1 port map( A => registers_1_22_port, ZN => n1319);
   U2165 : INV_X1 port map( A => registers_17_22_port, ZN => n1322);
   U2166 : INV_X1 port map( A => registers_3_22_port, ZN => n1329);
   U2167 : INV_X1 port map( A => registers_9_21_port, ZN => n1280);
   U2168 : INV_X1 port map( A => registers_8_21_port, ZN => n1283);
   U2169 : INV_X1 port map( A => registers_1_21_port, ZN => n1286);
   U2170 : INV_X1 port map( A => registers_17_21_port, ZN => n1289);
   U2171 : INV_X1 port map( A => registers_3_21_port, ZN => n1296);
   U2172 : INV_X1 port map( A => registers_9_20_port, ZN => n1247);
   U2173 : INV_X1 port map( A => registers_8_20_port, ZN => n1250);
   U2174 : INV_X1 port map( A => registers_1_20_port, ZN => n1253);
   U2175 : INV_X1 port map( A => registers_17_20_port, ZN => n1256);
   U2176 : INV_X1 port map( A => registers_3_20_port, ZN => n1263);
   U2177 : INV_X1 port map( A => registers_9_19_port, ZN => n1214);
   U2178 : INV_X1 port map( A => registers_8_19_port, ZN => n1217);
   U2179 : INV_X1 port map( A => registers_1_19_port, ZN => n1220);
   U2180 : INV_X1 port map( A => registers_17_19_port, ZN => n1223);
   U2181 : INV_X1 port map( A => registers_3_19_port, ZN => n1230);
   U2182 : INV_X1 port map( A => registers_9_18_port, ZN => n1181);
   U2183 : INV_X1 port map( A => registers_8_18_port, ZN => n1184);
   U2184 : INV_X1 port map( A => registers_1_18_port, ZN => n1187);
   U2185 : INV_X1 port map( A => registers_17_18_port, ZN => n1190);
   U2186 : INV_X1 port map( A => registers_3_18_port, ZN => n1197);
   U2187 : INV_X1 port map( A => registers_9_17_port, ZN => n1148);
   U2188 : INV_X1 port map( A => registers_8_17_port, ZN => n1151);
   U2189 : INV_X1 port map( A => registers_1_17_port, ZN => n1154);
   U2190 : INV_X1 port map( A => registers_17_17_port, ZN => n1157);
   U2191 : INV_X1 port map( A => registers_3_17_port, ZN => n1164);
   U2192 : INV_X1 port map( A => registers_9_16_port, ZN => n1115);
   U2193 : INV_X1 port map( A => registers_8_16_port, ZN => n1118);
   U2194 : INV_X1 port map( A => registers_1_16_port, ZN => n1121);
   U2195 : INV_X1 port map( A => registers_17_16_port, ZN => n1124);
   U2196 : INV_X1 port map( A => registers_3_16_port, ZN => n1131);
   U2197 : AND2_X1 port map( A1 => data_in_port_w(0), A2 => n5179, ZN => n2976)
                           ;
   U2198 : AND2_X1 port map( A1 => data_in_port_w(1), A2 => n5179, ZN => n2979)
                           ;
   U2199 : AND2_X1 port map( A1 => data_in_port_w(2), A2 => n5179, ZN => n2982)
                           ;
   U2200 : AND2_X1 port map( A1 => data_in_port_w(3), A2 => n5179, ZN => n2985)
                           ;
   U2201 : AND2_X1 port map( A1 => data_in_port_w(4), A2 => n5179, ZN => n2988)
                           ;
   U2202 : AND2_X1 port map( A1 => data_in_port_w(5), A2 => n5179, ZN => n2991)
                           ;
   U2203 : AND2_X1 port map( A1 => data_in_port_w(6), A2 => n5179, ZN => n2994)
                           ;
   U2204 : AND2_X1 port map( A1 => data_in_port_w(7), A2 => n5179, ZN => n2997)
                           ;
   U2205 : AND2_X1 port map( A1 => data_in_port_w(8), A2 => n5180, ZN => n3000)
                           ;
   U2206 : AND2_X1 port map( A1 => data_in_port_w(9), A2 => n5180, ZN => n3003)
                           ;
   U2207 : AND2_X1 port map( A1 => data_in_port_w(10), A2 => n5180, ZN => n3006
                           );
   U2208 : AND2_X1 port map( A1 => data_in_port_w(11), A2 => n5180, ZN => n3009
                           );
   U2209 : AND2_X1 port map( A1 => data_in_port_w(12), A2 => n5180, ZN => n3012
                           );
   U2210 : AND2_X1 port map( A1 => data_in_port_w(13), A2 => n5180, ZN => n3015
                           );
   U2211 : AND2_X1 port map( A1 => data_in_port_w(14), A2 => n5180, ZN => n3018
                           );
   U2212 : AND2_X1 port map( A1 => data_in_port_w(15), A2 => n5180, ZN => n3021
                           );
   U2213 : AND2_X1 port map( A1 => data_in_port_w(16), A2 => n5180, ZN => n3024
                           );
   U2214 : AND2_X1 port map( A1 => data_in_port_w(17), A2 => n5180, ZN => n3027
                           );
   U2215 : AND2_X1 port map( A1 => data_in_port_w(18), A2 => n5180, ZN => n3030
                           );
   U2216 : AND2_X1 port map( A1 => data_in_port_w(19), A2 => n5180, ZN => n3033
                           );
   U2217 : AND2_X1 port map( A1 => data_in_port_w(20), A2 => n5180, ZN => n3036
                           );
   U2218 : AND2_X1 port map( A1 => data_in_port_w(21), A2 => n5180, ZN => n3039
                           );
   U2219 : AND2_X1 port map( A1 => data_in_port_w(22), A2 => n5180, ZN => n3042
                           );
   U2220 : AND2_X1 port map( A1 => data_in_port_w(23), A2 => n5180, ZN => n3045
                           );
   U2221 : AND2_X1 port map( A1 => data_in_port_w(24), A2 => n5180, ZN => n3048
                           );
   U2222 : AND2_X1 port map( A1 => data_in_port_w(25), A2 => n5180, ZN => n3051
                           );
   U2223 : AND2_X1 port map( A1 => data_in_port_w(26), A2 => n5181, ZN => n3054
                           );
   U2224 : AND2_X1 port map( A1 => data_in_port_w(27), A2 => n5181, ZN => n3057
                           );
   U2225 : AND2_X1 port map( A1 => data_in_port_w(28), A2 => n5181, ZN => n3060
                           );
   U2226 : AND2_X1 port map( A1 => data_in_port_w(29), A2 => n5181, ZN => n3063
                           );
   U2227 : AND2_X1 port map( A1 => data_in_port_w(30), A2 => n5181, ZN => n3066
                           );
   U2228 : AND2_X1 port map( A1 => data_in_port_w(31), A2 => n5181, ZN => n3069
                           );
   U2229 : INV_X1 port map( A => reset, ZN => n5182);
   U2230 : INV_X1 port map( A => address_port_w(4), ZN => n539);
   U2231 : INV_X1 port map( A => address_port_w(3), ZN => n538);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity hazardUnit is

   port( RS_address, RT_address, RT_address_ID_EX : in std_logic_vector (4 
         downto 0);  MemRead_ID_EX, multi_cycle_operation : in std_logic;  
         enable_signal, sel1 : out std_logic);

end hazardUnit;

architecture SYN_Behavioral of hazardUnit is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13 : 
      std_logic;

begin
   enable_signal <= sel1_port;
   sel1 <= sel1_port;
   
   U8 : OAI33_X1 port map( A1 => n2, A2 => n3, A3 => n4, B1 => n5, B2 => n6, B3
                           => n7, ZN => n1);
   U9 : XOR2_X1 port map( A => RT_address_ID_EX(4), B => RS_address(4), Z => n7
                           );
   U10 : XOR2_X1 port map( A => RT_address_ID_EX(2), B => RS_address(2), Z => 
                           n6);
   U11 : NAND3_X1 port map( A1 => n8, A2 => n9, A3 => n10, ZN => n5);
   U12 : XOR2_X1 port map( A => RT_address_ID_EX(4), B => RT_address(4), Z => 
                           n4);
   U13 : XOR2_X1 port map( A => RT_address_ID_EX(3), B => RT_address(3), Z => 
                           n3);
   U14 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => n2);
   U1 : AOI21_X1 port map( B1 => MemRead_ID_EX, B2 => n1, A => 
                           multi_cycle_operation, ZN => sel1_port);
   U2 : XNOR2_X1 port map( A => RT_address_ID_EX(0), B => RT_address(0), ZN => 
                           n12);
   U3 : XNOR2_X1 port map( A => RT_address_ID_EX(0), B => RS_address(0), ZN => 
                           n9);
   U4 : XNOR2_X1 port map( A => RT_address_ID_EX(3), B => RS_address(3), ZN => 
                           n8);
   U5 : XNOR2_X1 port map( A => RT_address_ID_EX(1), B => RT_address(1), ZN => 
                           n13);
   U6 : XNOR2_X1 port map( A => RT_address_ID_EX(1), B => RS_address(1), ZN => 
                           n10);
   U7 : XNOR2_X1 port map( A => RT_address_ID_EX(2), B => RT_address(2), ZN => 
                           n11);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity comparator is

   port( A, B : in std_logic_vector (31 downto 0);  Sel : in std_logic_vector 
         (2 downto 0);  O : out std_logic_vector (31 downto 0));

end comparator;

architecture SYN_Behavioral of comparator is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator_DW01_cmp6_1
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component comparator_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_0_port, N14, N19, N20, net166336, net166335, 
      net166334, net166333, net166332, net166331, net166330, net166329, 
      net166328, n3, n4, n8, n9, n10, n11, n12, n13, n14_port, n15 : std_logic;

begin
   O <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, O_0_port );
   
   X_Logic0_port <= '0';
   n3 <= '1';
   n4 <= '0';
   U14 : NAND3_X1 port map( A1 => n10, A2 => n11, A3 => Sel(2), ZN => n9);
   r71 : comparator_DW01_cmp6_0 port map( A(31) => B(31), A(30) => B(30), A(29)
                           => B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B(31) => A(31), B(30) => A(30), B(29) => 
                           A(29), B(28) => A(28), B(27) => A(27), B(26) => 
                           A(26), B(25) => A(25), B(24) => A(24), B(23) => 
                           A(23), B(22) => A(22), B(21) => A(21), B(20) => 
                           A(20), B(19) => A(19), B(18) => A(18), B(17) => 
                           A(17), B(16) => A(16), B(15) => A(15), B(14) => 
                           A(14), B(13) => A(13), B(12) => A(12), B(11) => 
                           A(11), B(10) => A(10), B(9) => A(9), B(8) => A(8), 
                           B(7) => A(7), B(6) => A(6), B(5) => A(5), B(4) => 
                           A(4), B(3) => A(3), B(2) => A(2), B(1) => A(1), B(0)
                           => A(0), TC => n3, LT => net166333, GT => N19, EQ =>
                           net166334, LE => net166335, GE => N20, NE => 
                           net166336);
   r70 : comparator_DW01_cmp6_1 port map( A(31) => A(31), A(30) => A(30), A(29)
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), TC => n4, LT => net166328, GT => net166329,
                           EQ => N14, LE => net166330, GE => net166331, NE => 
                           net166332);
   U4 : INV_X1 port map( A => Sel(0), ZN => n13);
   U5 : OAI22_X1 port map( A1 => Sel(0), A2 => N20, B1 => N19, B2 => n13, ZN =>
                           n15);
   U6 : AOI22_X1 port map( A1 => n14_port, A2 => n11, B1 => Sel(1), B2 => n15, 
                           ZN => n8);
   U7 : INV_X1 port map( A => Sel(1), ZN => n11);
   U8 : XNOR2_X1 port map( A => n13, B => N14, ZN => n14_port);
   U9 : INV_X1 port map( A => n12, ZN => n10);
   U10 : AOI22_X1 port map( A1 => N20, A2 => Sel(0), B1 => n13, B2 => N19, ZN 
                           => n12);
   U11 : OAI21_X1 port map( B1 => Sel(2), B2 => n8, A => n9, ZN => O_0_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity logicUnitT2_data_size32 is

   port( operand_a, operand_b : in std_logic_vector (31 downto 0);  type_op : 
         in std_logic_vector (3 downto 0);  result : out std_logic_vector (31 
         downto 0));

end logicUnitT2_data_size32;

architecture SYN_Behavioral of logicUnitT2_data_size32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component nandWithEn_data_size32_1
      port( operand_a, operand_b : in std_logic_vector (31 downto 0);  enable :
            in std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component nandWithEn_data_size32_2
      port( operand_a, operand_b : in std_logic_vector (31 downto 0);  enable :
            in std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component nandWithEn_data_size32_3
      port( operand_a, operand_b : in std_logic_vector (31 downto 0);  enable :
            in std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component nandWithEn_data_size32_0
      port( operand_a, operand_b : in std_logic_vector (31 downto 0);  enable :
            in std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   signal notA_31_port, notA_30_port, notA_29_port, notA_28_port, notA_27_port,
      notA_26_port, notA_25_port, notA_24_port, notA_23_port, notA_22_port, 
      notA_21_port, notA_20_port, notA_19_port, notA_18_port, notA_17_port, 
      notA_16_port, notA_15_port, notA_14_port, notA_13_port, notA_12_port, 
      notA_11_port, notA_10_port, notA_9_port, notA_8_port, notA_7_port, 
      notA_6_port, notA_5_port, notA_4_port, notA_3_port, notA_2_port, 
      notA_1_port, notA_0_port, notB_31_port, notB_30_port, notB_29_port, 
      notB_28_port, notB_27_port, notB_26_port, notB_25_port, notB_24_port, 
      notB_23_port, notB_22_port, notB_21_port, notB_20_port, notB_19_port, 
      notB_18_port, notB_17_port, notB_16_port, notB_15_port, notB_14_port, 
      notB_13_port, notB_12_port, notB_11_port, notB_10_port, notB_9_port, 
      notB_8_port, notB_7_port, notB_6_port, notB_5_port, notB_4_port, 
      notB_3_port, notB_2_port, notB_1_port, notB_0_port, 
      partial_result_l0_31_port, partial_result_l0_30_port, 
      partial_result_l0_29_port, partial_result_l0_28_port, 
      partial_result_l0_27_port, partial_result_l0_26_port, 
      partial_result_l0_25_port, partial_result_l0_24_port, 
      partial_result_l0_23_port, partial_result_l0_22_port, 
      partial_result_l0_21_port, partial_result_l0_20_port, 
      partial_result_l0_19_port, partial_result_l0_18_port, 
      partial_result_l0_17_port, partial_result_l0_16_port, 
      partial_result_l0_15_port, partial_result_l0_14_port, 
      partial_result_l0_13_port, partial_result_l0_12_port, 
      partial_result_l0_11_port, partial_result_l0_10_port, 
      partial_result_l0_9_port, partial_result_l0_8_port, 
      partial_result_l0_7_port, partial_result_l0_6_port, 
      partial_result_l0_5_port, partial_result_l0_4_port, 
      partial_result_l0_3_port, partial_result_l0_2_port, 
      partial_result_l0_1_port, partial_result_l0_0_port, 
      partial_result_l1_31_port, partial_result_l1_30_port, 
      partial_result_l1_29_port, partial_result_l1_28_port, 
      partial_result_l1_27_port, partial_result_l1_26_port, 
      partial_result_l1_25_port, partial_result_l1_24_port, 
      partial_result_l1_23_port, partial_result_l1_22_port, 
      partial_result_l1_21_port, partial_result_l1_20_port, 
      partial_result_l1_19_port, partial_result_l1_18_port, 
      partial_result_l1_17_port, partial_result_l1_16_port, 
      partial_result_l1_15_port, partial_result_l1_14_port, 
      partial_result_l1_13_port, partial_result_l1_12_port, 
      partial_result_l1_11_port, partial_result_l1_10_port, 
      partial_result_l1_9_port, partial_result_l1_8_port, 
      partial_result_l1_7_port, partial_result_l1_6_port, 
      partial_result_l1_5_port, partial_result_l1_4_port, 
      partial_result_l1_3_port, partial_result_l1_2_port, 
      partial_result_l1_1_port, partial_result_l1_0_port, 
      partial_result_l2_31_port, partial_result_l2_30_port, 
      partial_result_l2_29_port, partial_result_l2_28_port, 
      partial_result_l2_27_port, partial_result_l2_26_port, 
      partial_result_l2_25_port, partial_result_l2_24_port, 
      partial_result_l2_23_port, partial_result_l2_22_port, 
      partial_result_l2_21_port, partial_result_l2_20_port, 
      partial_result_l2_19_port, partial_result_l2_18_port, 
      partial_result_l2_17_port, partial_result_l2_16_port, 
      partial_result_l2_15_port, partial_result_l2_14_port, 
      partial_result_l2_13_port, partial_result_l2_12_port, 
      partial_result_l2_11_port, partial_result_l2_10_port, 
      partial_result_l2_9_port, partial_result_l2_8_port, 
      partial_result_l2_7_port, partial_result_l2_6_port, 
      partial_result_l2_5_port, partial_result_l2_4_port, 
      partial_result_l2_3_port, partial_result_l2_2_port, 
      partial_result_l2_1_port, partial_result_l2_0_port, 
      partial_result_l3_31_port, partial_result_l3_30_port, 
      partial_result_l3_29_port, partial_result_l3_28_port, 
      partial_result_l3_27_port, partial_result_l3_26_port, 
      partial_result_l3_25_port, partial_result_l3_24_port, 
      partial_result_l3_23_port, partial_result_l3_22_port, 
      partial_result_l3_21_port, partial_result_l3_20_port, 
      partial_result_l3_19_port, partial_result_l3_18_port, 
      partial_result_l3_17_port, partial_result_l3_16_port, 
      partial_result_l3_15_port, partial_result_l3_14_port, 
      partial_result_l3_13_port, partial_result_l3_12_port, 
      partial_result_l3_11_port, partial_result_l3_10_port, 
      partial_result_l3_9_port, partial_result_l3_8_port, 
      partial_result_l3_7_port, partial_result_l3_6_port, 
      partial_result_l3_5_port, partial_result_l3_4_port, 
      partial_result_l3_3_port, partial_result_l3_2_port, 
      partial_result_l3_1_port, partial_result_l3_0_port : std_logic;

begin
   
   n0 : nandWithEn_data_size32_0 port map( operand_a(31) => notA_31_port, 
                           operand_a(30) => notA_30_port, operand_a(29) => 
                           notA_29_port, operand_a(28) => notA_28_port, 
                           operand_a(27) => notA_27_port, operand_a(26) => 
                           notA_26_port, operand_a(25) => notA_25_port, 
                           operand_a(24) => notA_24_port, operand_a(23) => 
                           notA_23_port, operand_a(22) => notA_22_port, 
                           operand_a(21) => notA_21_port, operand_a(20) => 
                           notA_20_port, operand_a(19) => notA_19_port, 
                           operand_a(18) => notA_18_port, operand_a(17) => 
                           notA_17_port, operand_a(16) => notA_16_port, 
                           operand_a(15) => notA_15_port, operand_a(14) => 
                           notA_14_port, operand_a(13) => notA_13_port, 
                           operand_a(12) => notA_12_port, operand_a(11) => 
                           notA_11_port, operand_a(10) => notA_10_port, 
                           operand_a(9) => notA_9_port, operand_a(8) => 
                           notA_8_port, operand_a(7) => notA_7_port, 
                           operand_a(6) => notA_6_port, operand_a(5) => 
                           notA_5_port, operand_a(4) => notA_4_port, 
                           operand_a(3) => notA_3_port, operand_a(2) => 
                           notA_2_port, operand_a(1) => notA_1_port, 
                           operand_a(0) => notA_0_port, operand_b(31) => 
                           notB_31_port, operand_b(30) => notB_30_port, 
                           operand_b(29) => notB_29_port, operand_b(28) => 
                           notB_28_port, operand_b(27) => notB_27_port, 
                           operand_b(26) => notB_26_port, operand_b(25) => 
                           notB_25_port, operand_b(24) => notB_24_port, 
                           operand_b(23) => notB_23_port, operand_b(22) => 
                           notB_22_port, operand_b(21) => notB_21_port, 
                           operand_b(20) => notB_20_port, operand_b(19) => 
                           notB_19_port, operand_b(18) => notB_18_port, 
                           operand_b(17) => notB_17_port, operand_b(16) => 
                           notB_16_port, operand_b(15) => notB_15_port, 
                           operand_b(14) => notB_14_port, operand_b(13) => 
                           notB_13_port, operand_b(12) => notB_12_port, 
                           operand_b(11) => notB_11_port, operand_b(10) => 
                           notB_10_port, operand_b(9) => notB_9_port, 
                           operand_b(8) => notB_8_port, operand_b(7) => 
                           notB_7_port, operand_b(6) => notB_6_port, 
                           operand_b(5) => notB_5_port, operand_b(4) => 
                           notB_4_port, operand_b(3) => notB_3_port, 
                           operand_b(2) => notB_2_port, operand_b(1) => 
                           notB_1_port, operand_b(0) => notB_0_port, enable => 
                           type_op(0), output(31) => partial_result_l0_31_port,
                           output(30) => partial_result_l0_30_port, output(29) 
                           => partial_result_l0_29_port, output(28) => 
                           partial_result_l0_28_port, output(27) => 
                           partial_result_l0_27_port, output(26) => 
                           partial_result_l0_26_port, output(25) => 
                           partial_result_l0_25_port, output(24) => 
                           partial_result_l0_24_port, output(23) => 
                           partial_result_l0_23_port, output(22) => 
                           partial_result_l0_22_port, output(21) => 
                           partial_result_l0_21_port, output(20) => 
                           partial_result_l0_20_port, output(19) => 
                           partial_result_l0_19_port, output(18) => 
                           partial_result_l0_18_port, output(17) => 
                           partial_result_l0_17_port, output(16) => 
                           partial_result_l0_16_port, output(15) => 
                           partial_result_l0_15_port, output(14) => 
                           partial_result_l0_14_port, output(13) => 
                           partial_result_l0_13_port, output(12) => 
                           partial_result_l0_12_port, output(11) => 
                           partial_result_l0_11_port, output(10) => 
                           partial_result_l0_10_port, output(9) => 
                           partial_result_l0_9_port, output(8) => 
                           partial_result_l0_8_port, output(7) => 
                           partial_result_l0_7_port, output(6) => 
                           partial_result_l0_6_port, output(5) => 
                           partial_result_l0_5_port, output(4) => 
                           partial_result_l0_4_port, output(3) => 
                           partial_result_l0_3_port, output(2) => 
                           partial_result_l0_2_port, output(1) => 
                           partial_result_l0_1_port, output(0) => 
                           partial_result_l0_0_port);
   n1 : nandWithEn_data_size32_3 port map( operand_a(31) => operand_a(31), 
                           operand_a(30) => operand_a(30), operand_a(29) => 
                           operand_a(29), operand_a(28) => operand_a(28), 
                           operand_a(27) => operand_a(27), operand_a(26) => 
                           operand_a(26), operand_a(25) => operand_a(25), 
                           operand_a(24) => operand_a(24), operand_a(23) => 
                           operand_a(23), operand_a(22) => operand_a(22), 
                           operand_a(21) => operand_a(21), operand_a(20) => 
                           operand_a(20), operand_a(19) => operand_a(19), 
                           operand_a(18) => operand_a(18), operand_a(17) => 
                           operand_a(17), operand_a(16) => operand_a(16), 
                           operand_a(15) => operand_a(15), operand_a(14) => 
                           operand_a(14), operand_a(13) => operand_a(13), 
                           operand_a(12) => operand_a(12), operand_a(11) => 
                           operand_a(11), operand_a(10) => operand_a(10), 
                           operand_a(9) => operand_a(9), operand_a(8) => 
                           operand_a(8), operand_a(7) => operand_a(7), 
                           operand_a(6) => operand_a(6), operand_a(5) => 
                           operand_a(5), operand_a(4) => operand_a(4), 
                           operand_a(3) => operand_a(3), operand_a(2) => 
                           operand_a(2), operand_a(1) => operand_a(1), 
                           operand_a(0) => operand_a(0), operand_b(31) => 
                           notB_31_port, operand_b(30) => notB_30_port, 
                           operand_b(29) => notB_29_port, operand_b(28) => 
                           notB_28_port, operand_b(27) => notB_27_port, 
                           operand_b(26) => notB_26_port, operand_b(25) => 
                           notB_25_port, operand_b(24) => notB_24_port, 
                           operand_b(23) => notB_23_port, operand_b(22) => 
                           notB_22_port, operand_b(21) => notB_21_port, 
                           operand_b(20) => notB_20_port, operand_b(19) => 
                           notB_19_port, operand_b(18) => notB_18_port, 
                           operand_b(17) => notB_17_port, operand_b(16) => 
                           notB_16_port, operand_b(15) => notB_15_port, 
                           operand_b(14) => notB_14_port, operand_b(13) => 
                           notB_13_port, operand_b(12) => notB_12_port, 
                           operand_b(11) => notB_11_port, operand_b(10) => 
                           notB_10_port, operand_b(9) => notB_9_port, 
                           operand_b(8) => notB_8_port, operand_b(7) => 
                           notB_7_port, operand_b(6) => notB_6_port, 
                           operand_b(5) => notB_5_port, operand_b(4) => 
                           notB_4_port, operand_b(3) => notB_3_port, 
                           operand_b(2) => notB_2_port, operand_b(1) => 
                           notB_1_port, operand_b(0) => notB_0_port, enable => 
                           type_op(1), output(31) => partial_result_l1_31_port,
                           output(30) => partial_result_l1_30_port, output(29) 
                           => partial_result_l1_29_port, output(28) => 
                           partial_result_l1_28_port, output(27) => 
                           partial_result_l1_27_port, output(26) => 
                           partial_result_l1_26_port, output(25) => 
                           partial_result_l1_25_port, output(24) => 
                           partial_result_l1_24_port, output(23) => 
                           partial_result_l1_23_port, output(22) => 
                           partial_result_l1_22_port, output(21) => 
                           partial_result_l1_21_port, output(20) => 
                           partial_result_l1_20_port, output(19) => 
                           partial_result_l1_19_port, output(18) => 
                           partial_result_l1_18_port, output(17) => 
                           partial_result_l1_17_port, output(16) => 
                           partial_result_l1_16_port, output(15) => 
                           partial_result_l1_15_port, output(14) => 
                           partial_result_l1_14_port, output(13) => 
                           partial_result_l1_13_port, output(12) => 
                           partial_result_l1_12_port, output(11) => 
                           partial_result_l1_11_port, output(10) => 
                           partial_result_l1_10_port, output(9) => 
                           partial_result_l1_9_port, output(8) => 
                           partial_result_l1_8_port, output(7) => 
                           partial_result_l1_7_port, output(6) => 
                           partial_result_l1_6_port, output(5) => 
                           partial_result_l1_5_port, output(4) => 
                           partial_result_l1_4_port, output(3) => 
                           partial_result_l1_3_port, output(2) => 
                           partial_result_l1_2_port, output(1) => 
                           partial_result_l1_1_port, output(0) => 
                           partial_result_l1_0_port);
   n2 : nandWithEn_data_size32_2 port map( operand_a(31) => notA_31_port, 
                           operand_a(30) => notA_30_port, operand_a(29) => 
                           notA_29_port, operand_a(28) => notA_28_port, 
                           operand_a(27) => notA_27_port, operand_a(26) => 
                           notA_26_port, operand_a(25) => notA_25_port, 
                           operand_a(24) => notA_24_port, operand_a(23) => 
                           notA_23_port, operand_a(22) => notA_22_port, 
                           operand_a(21) => notA_21_port, operand_a(20) => 
                           notA_20_port, operand_a(19) => notA_19_port, 
                           operand_a(18) => notA_18_port, operand_a(17) => 
                           notA_17_port, operand_a(16) => notA_16_port, 
                           operand_a(15) => notA_15_port, operand_a(14) => 
                           notA_14_port, operand_a(13) => notA_13_port, 
                           operand_a(12) => notA_12_port, operand_a(11) => 
                           notA_11_port, operand_a(10) => notA_10_port, 
                           operand_a(9) => notA_9_port, operand_a(8) => 
                           notA_8_port, operand_a(7) => notA_7_port, 
                           operand_a(6) => notA_6_port, operand_a(5) => 
                           notA_5_port, operand_a(4) => notA_4_port, 
                           operand_a(3) => notA_3_port, operand_a(2) => 
                           notA_2_port, operand_a(1) => notA_1_port, 
                           operand_a(0) => notA_0_port, operand_b(31) => 
                           operand_b(31), operand_b(30) => operand_b(30), 
                           operand_b(29) => operand_b(29), operand_b(28) => 
                           operand_b(28), operand_b(27) => operand_b(27), 
                           operand_b(26) => operand_b(26), operand_b(25) => 
                           operand_b(25), operand_b(24) => operand_b(24), 
                           operand_b(23) => operand_b(23), operand_b(22) => 
                           operand_b(22), operand_b(21) => operand_b(21), 
                           operand_b(20) => operand_b(20), operand_b(19) => 
                           operand_b(19), operand_b(18) => operand_b(18), 
                           operand_b(17) => operand_b(17), operand_b(16) => 
                           operand_b(16), operand_b(15) => operand_b(15), 
                           operand_b(14) => operand_b(14), operand_b(13) => 
                           operand_b(13), operand_b(12) => operand_b(12), 
                           operand_b(11) => operand_b(11), operand_b(10) => 
                           operand_b(10), operand_b(9) => operand_b(9), 
                           operand_b(8) => operand_b(8), operand_b(7) => 
                           operand_b(7), operand_b(6) => operand_b(6), 
                           operand_b(5) => operand_b(5), operand_b(4) => 
                           operand_b(4), operand_b(3) => operand_b(3), 
                           operand_b(2) => operand_b(2), operand_b(1) => 
                           operand_b(1), operand_b(0) => operand_b(0), enable 
                           => type_op(2), output(31) => 
                           partial_result_l2_31_port, output(30) => 
                           partial_result_l2_30_port, output(29) => 
                           partial_result_l2_29_port, output(28) => 
                           partial_result_l2_28_port, output(27) => 
                           partial_result_l2_27_port, output(26) => 
                           partial_result_l2_26_port, output(25) => 
                           partial_result_l2_25_port, output(24) => 
                           partial_result_l2_24_port, output(23) => 
                           partial_result_l2_23_port, output(22) => 
                           partial_result_l2_22_port, output(21) => 
                           partial_result_l2_21_port, output(20) => 
                           partial_result_l2_20_port, output(19) => 
                           partial_result_l2_19_port, output(18) => 
                           partial_result_l2_18_port, output(17) => 
                           partial_result_l2_17_port, output(16) => 
                           partial_result_l2_16_port, output(15) => 
                           partial_result_l2_15_port, output(14) => 
                           partial_result_l2_14_port, output(13) => 
                           partial_result_l2_13_port, output(12) => 
                           partial_result_l2_12_port, output(11) => 
                           partial_result_l2_11_port, output(10) => 
                           partial_result_l2_10_port, output(9) => 
                           partial_result_l2_9_port, output(8) => 
                           partial_result_l2_8_port, output(7) => 
                           partial_result_l2_7_port, output(6) => 
                           partial_result_l2_6_port, output(5) => 
                           partial_result_l2_5_port, output(4) => 
                           partial_result_l2_4_port, output(3) => 
                           partial_result_l2_3_port, output(2) => 
                           partial_result_l2_2_port, output(1) => 
                           partial_result_l2_1_port, output(0) => 
                           partial_result_l2_0_port);
   n3 : nandWithEn_data_size32_1 port map( operand_a(31) => operand_a(31), 
                           operand_a(30) => operand_a(30), operand_a(29) => 
                           operand_a(29), operand_a(28) => operand_a(28), 
                           operand_a(27) => operand_a(27), operand_a(26) => 
                           operand_a(26), operand_a(25) => operand_a(25), 
                           operand_a(24) => operand_a(24), operand_a(23) => 
                           operand_a(23), operand_a(22) => operand_a(22), 
                           operand_a(21) => operand_a(21), operand_a(20) => 
                           operand_a(20), operand_a(19) => operand_a(19), 
                           operand_a(18) => operand_a(18), operand_a(17) => 
                           operand_a(17), operand_a(16) => operand_a(16), 
                           operand_a(15) => operand_a(15), operand_a(14) => 
                           operand_a(14), operand_a(13) => operand_a(13), 
                           operand_a(12) => operand_a(12), operand_a(11) => 
                           operand_a(11), operand_a(10) => operand_a(10), 
                           operand_a(9) => operand_a(9), operand_a(8) => 
                           operand_a(8), operand_a(7) => operand_a(7), 
                           operand_a(6) => operand_a(6), operand_a(5) => 
                           operand_a(5), operand_a(4) => operand_a(4), 
                           operand_a(3) => operand_a(3), operand_a(2) => 
                           operand_a(2), operand_a(1) => operand_a(1), 
                           operand_a(0) => operand_a(0), operand_b(31) => 
                           operand_b(31), operand_b(30) => operand_b(30), 
                           operand_b(29) => operand_b(29), operand_b(28) => 
                           operand_b(28), operand_b(27) => operand_b(27), 
                           operand_b(26) => operand_b(26), operand_b(25) => 
                           operand_b(25), operand_b(24) => operand_b(24), 
                           operand_b(23) => operand_b(23), operand_b(22) => 
                           operand_b(22), operand_b(21) => operand_b(21), 
                           operand_b(20) => operand_b(20), operand_b(19) => 
                           operand_b(19), operand_b(18) => operand_b(18), 
                           operand_b(17) => operand_b(17), operand_b(16) => 
                           operand_b(16), operand_b(15) => operand_b(15), 
                           operand_b(14) => operand_b(14), operand_b(13) => 
                           operand_b(13), operand_b(12) => operand_b(12), 
                           operand_b(11) => operand_b(11), operand_b(10) => 
                           operand_b(10), operand_b(9) => operand_b(9), 
                           operand_b(8) => operand_b(8), operand_b(7) => 
                           operand_b(7), operand_b(6) => operand_b(6), 
                           operand_b(5) => operand_b(5), operand_b(4) => 
                           operand_b(4), operand_b(3) => operand_b(3), 
                           operand_b(2) => operand_b(2), operand_b(1) => 
                           operand_b(1), operand_b(0) => operand_b(0), enable 
                           => type_op(3), output(31) => 
                           partial_result_l3_31_port, output(30) => 
                           partial_result_l3_30_port, output(29) => 
                           partial_result_l3_29_port, output(28) => 
                           partial_result_l3_28_port, output(27) => 
                           partial_result_l3_27_port, output(26) => 
                           partial_result_l3_26_port, output(25) => 
                           partial_result_l3_25_port, output(24) => 
                           partial_result_l3_24_port, output(23) => 
                           partial_result_l3_23_port, output(22) => 
                           partial_result_l3_22_port, output(21) => 
                           partial_result_l3_21_port, output(20) => 
                           partial_result_l3_20_port, output(19) => 
                           partial_result_l3_19_port, output(18) => 
                           partial_result_l3_18_port, output(17) => 
                           partial_result_l3_17_port, output(16) => 
                           partial_result_l3_16_port, output(15) => 
                           partial_result_l3_15_port, output(14) => 
                           partial_result_l3_14_port, output(13) => 
                           partial_result_l3_13_port, output(12) => 
                           partial_result_l3_12_port, output(11) => 
                           partial_result_l3_11_port, output(10) => 
                           partial_result_l3_10_port, output(9) => 
                           partial_result_l3_9_port, output(8) => 
                           partial_result_l3_8_port, output(7) => 
                           partial_result_l3_7_port, output(6) => 
                           partial_result_l3_6_port, output(5) => 
                           partial_result_l3_5_port, output(4) => 
                           partial_result_l3_4_port, output(3) => 
                           partial_result_l3_3_port, output(2) => 
                           partial_result_l3_2_port, output(1) => 
                           partial_result_l3_1_port, output(0) => 
                           partial_result_l3_0_port);
   U1 : NAND4_X1 port map( A1 => partial_result_l3_15_port, A2 => 
                           partial_result_l2_15_port, A3 => 
                           partial_result_l1_15_port, A4 => 
                           partial_result_l0_15_port, ZN => result(15));
   U2 : NAND4_X1 port map( A1 => partial_result_l3_14_port, A2 => 
                           partial_result_l2_14_port, A3 => 
                           partial_result_l1_14_port, A4 => 
                           partial_result_l0_14_port, ZN => result(14));
   U3 : NAND4_X1 port map( A1 => partial_result_l3_13_port, A2 => 
                           partial_result_l2_13_port, A3 => 
                           partial_result_l1_13_port, A4 => 
                           partial_result_l0_13_port, ZN => result(13));
   U4 : NAND4_X1 port map( A1 => partial_result_l3_12_port, A2 => 
                           partial_result_l2_12_port, A3 => 
                           partial_result_l1_12_port, A4 => 
                           partial_result_l0_12_port, ZN => result(12));
   U5 : NAND4_X1 port map( A1 => partial_result_l3_11_port, A2 => 
                           partial_result_l2_11_port, A3 => 
                           partial_result_l1_11_port, A4 => 
                           partial_result_l0_11_port, ZN => result(11));
   U6 : NAND4_X1 port map( A1 => partial_result_l3_10_port, A2 => 
                           partial_result_l2_10_port, A3 => 
                           partial_result_l1_10_port, A4 => 
                           partial_result_l0_10_port, ZN => result(10));
   U7 : NAND4_X1 port map( A1 => partial_result_l3_9_port, A2 => 
                           partial_result_l2_9_port, A3 => 
                           partial_result_l1_9_port, A4 => 
                           partial_result_l0_9_port, ZN => result(9));
   U8 : NAND4_X1 port map( A1 => partial_result_l3_8_port, A2 => 
                           partial_result_l2_8_port, A3 => 
                           partial_result_l1_8_port, A4 => 
                           partial_result_l0_8_port, ZN => result(8));
   U9 : NAND4_X1 port map( A1 => partial_result_l3_7_port, A2 => 
                           partial_result_l2_7_port, A3 => 
                           partial_result_l1_7_port, A4 => 
                           partial_result_l0_7_port, ZN => result(7));
   U10 : NAND4_X1 port map( A1 => partial_result_l3_6_port, A2 => 
                           partial_result_l2_6_port, A3 => 
                           partial_result_l1_6_port, A4 => 
                           partial_result_l0_6_port, ZN => result(6));
   U11 : NAND4_X1 port map( A1 => partial_result_l3_5_port, A2 => 
                           partial_result_l2_5_port, A3 => 
                           partial_result_l1_5_port, A4 => 
                           partial_result_l0_5_port, ZN => result(5));
   U12 : NAND4_X1 port map( A1 => partial_result_l3_4_port, A2 => 
                           partial_result_l2_4_port, A3 => 
                           partial_result_l1_4_port, A4 => 
                           partial_result_l0_4_port, ZN => result(4));
   U13 : NAND4_X1 port map( A1 => partial_result_l3_3_port, A2 => 
                           partial_result_l2_3_port, A3 => 
                           partial_result_l1_3_port, A4 => 
                           partial_result_l0_3_port, ZN => result(3));
   U14 : NAND4_X1 port map( A1 => partial_result_l3_2_port, A2 => 
                           partial_result_l2_2_port, A3 => 
                           partial_result_l1_2_port, A4 => 
                           partial_result_l0_2_port, ZN => result(2));
   U15 : NAND4_X1 port map( A1 => partial_result_l3_1_port, A2 => 
                           partial_result_l2_1_port, A3 => 
                           partial_result_l1_1_port, A4 => 
                           partial_result_l0_1_port, ZN => result(1));
   U16 : NAND4_X1 port map( A1 => partial_result_l3_0_port, A2 => 
                           partial_result_l2_0_port, A3 => 
                           partial_result_l1_0_port, A4 => 
                           partial_result_l0_0_port, ZN => result(0));
   U17 : NAND4_X1 port map( A1 => partial_result_l3_31_port, A2 => 
                           partial_result_l2_31_port, A3 => 
                           partial_result_l1_31_port, A4 => 
                           partial_result_l0_31_port, ZN => result(31));
   U18 : NAND4_X1 port map( A1 => partial_result_l3_30_port, A2 => 
                           partial_result_l2_30_port, A3 => 
                           partial_result_l1_30_port, A4 => 
                           partial_result_l0_30_port, ZN => result(30));
   U19 : NAND4_X1 port map( A1 => partial_result_l3_29_port, A2 => 
                           partial_result_l2_29_port, A3 => 
                           partial_result_l1_29_port, A4 => 
                           partial_result_l0_29_port, ZN => result(29));
   U20 : NAND4_X1 port map( A1 => partial_result_l3_28_port, A2 => 
                           partial_result_l2_28_port, A3 => 
                           partial_result_l1_28_port, A4 => 
                           partial_result_l0_28_port, ZN => result(28));
   U21 : NAND4_X1 port map( A1 => partial_result_l3_27_port, A2 => 
                           partial_result_l2_27_port, A3 => 
                           partial_result_l1_27_port, A4 => 
                           partial_result_l0_27_port, ZN => result(27));
   U22 : NAND4_X1 port map( A1 => partial_result_l3_26_port, A2 => 
                           partial_result_l2_26_port, A3 => 
                           partial_result_l1_26_port, A4 => 
                           partial_result_l0_26_port, ZN => result(26));
   U23 : NAND4_X1 port map( A1 => partial_result_l3_25_port, A2 => 
                           partial_result_l2_25_port, A3 => 
                           partial_result_l1_25_port, A4 => 
                           partial_result_l0_25_port, ZN => result(25));
   U24 : NAND4_X1 port map( A1 => partial_result_l3_24_port, A2 => 
                           partial_result_l2_24_port, A3 => 
                           partial_result_l1_24_port, A4 => 
                           partial_result_l0_24_port, ZN => result(24));
   U25 : NAND4_X1 port map( A1 => partial_result_l3_23_port, A2 => 
                           partial_result_l2_23_port, A3 => 
                           partial_result_l1_23_port, A4 => 
                           partial_result_l0_23_port, ZN => result(23));
   U26 : NAND4_X1 port map( A1 => partial_result_l3_22_port, A2 => 
                           partial_result_l2_22_port, A3 => 
                           partial_result_l1_22_port, A4 => 
                           partial_result_l0_22_port, ZN => result(22));
   U27 : NAND4_X1 port map( A1 => partial_result_l3_21_port, A2 => 
                           partial_result_l2_21_port, A3 => 
                           partial_result_l1_21_port, A4 => 
                           partial_result_l0_21_port, ZN => result(21));
   U28 : NAND4_X1 port map( A1 => partial_result_l3_20_port, A2 => 
                           partial_result_l2_20_port, A3 => 
                           partial_result_l1_20_port, A4 => 
                           partial_result_l0_20_port, ZN => result(20));
   U29 : NAND4_X1 port map( A1 => partial_result_l3_19_port, A2 => 
                           partial_result_l2_19_port, A3 => 
                           partial_result_l1_19_port, A4 => 
                           partial_result_l0_19_port, ZN => result(19));
   U30 : NAND4_X1 port map( A1 => partial_result_l3_18_port, A2 => 
                           partial_result_l2_18_port, A3 => 
                           partial_result_l1_18_port, A4 => 
                           partial_result_l0_18_port, ZN => result(18));
   U31 : NAND4_X1 port map( A1 => partial_result_l3_17_port, A2 => 
                           partial_result_l2_17_port, A3 => 
                           partial_result_l1_17_port, A4 => 
                           partial_result_l0_17_port, ZN => result(17));
   U32 : NAND4_X1 port map( A1 => partial_result_l3_16_port, A2 => 
                           partial_result_l2_16_port, A3 => 
                           partial_result_l1_16_port, A4 => 
                           partial_result_l0_16_port, ZN => result(16));
   U33 : INV_X1 port map( A => operand_b(0), ZN => notB_0_port);
   U34 : INV_X1 port map( A => operand_b(1), ZN => notB_1_port);
   U35 : INV_X1 port map( A => operand_b(2), ZN => notB_2_port);
   U36 : INV_X1 port map( A => operand_b(3), ZN => notB_3_port);
   U37 : INV_X1 port map( A => operand_b(4), ZN => notB_4_port);
   U38 : INV_X1 port map( A => operand_b(5), ZN => notB_5_port);
   U39 : INV_X1 port map( A => operand_b(6), ZN => notB_6_port);
   U40 : INV_X1 port map( A => operand_b(7), ZN => notB_7_port);
   U41 : INV_X1 port map( A => operand_b(8), ZN => notB_8_port);
   U42 : INV_X1 port map( A => operand_b(9), ZN => notB_9_port);
   U43 : INV_X1 port map( A => operand_b(10), ZN => notB_10_port);
   U44 : INV_X1 port map( A => operand_b(11), ZN => notB_11_port);
   U45 : INV_X1 port map( A => operand_b(12), ZN => notB_12_port);
   U46 : INV_X1 port map( A => operand_b(13), ZN => notB_13_port);
   U47 : INV_X1 port map( A => operand_b(14), ZN => notB_14_port);
   U48 : INV_X1 port map( A => operand_b(15), ZN => notB_15_port);
   U49 : INV_X1 port map( A => operand_b(16), ZN => notB_16_port);
   U50 : INV_X1 port map( A => operand_b(17), ZN => notB_17_port);
   U51 : INV_X1 port map( A => operand_b(18), ZN => notB_18_port);
   U52 : INV_X1 port map( A => operand_b(19), ZN => notB_19_port);
   U53 : INV_X1 port map( A => operand_b(20), ZN => notB_20_port);
   U54 : INV_X1 port map( A => operand_b(21), ZN => notB_21_port);
   U55 : INV_X1 port map( A => operand_b(22), ZN => notB_22_port);
   U56 : INV_X1 port map( A => operand_b(23), ZN => notB_23_port);
   U57 : INV_X1 port map( A => operand_b(24), ZN => notB_24_port);
   U58 : INV_X1 port map( A => operand_b(25), ZN => notB_25_port);
   U59 : INV_X1 port map( A => operand_b(26), ZN => notB_26_port);
   U60 : INV_X1 port map( A => operand_b(27), ZN => notB_27_port);
   U61 : INV_X1 port map( A => operand_b(28), ZN => notB_28_port);
   U62 : INV_X1 port map( A => operand_b(29), ZN => notB_29_port);
   U63 : INV_X1 port map( A => operand_b(30), ZN => notB_30_port);
   U64 : INV_X1 port map( A => operand_b(31), ZN => notB_31_port);
   U65 : INV_X1 port map( A => operand_a(0), ZN => notA_0_port);
   U66 : INV_X1 port map( A => operand_a(1), ZN => notA_1_port);
   U67 : INV_X1 port map( A => operand_a(2), ZN => notA_2_port);
   U68 : INV_X1 port map( A => operand_a(3), ZN => notA_3_port);
   U69 : INV_X1 port map( A => operand_a(4), ZN => notA_4_port);
   U70 : INV_X1 port map( A => operand_a(5), ZN => notA_5_port);
   U71 : INV_X1 port map( A => operand_a(6), ZN => notA_6_port);
   U72 : INV_X1 port map( A => operand_a(7), ZN => notA_7_port);
   U73 : INV_X1 port map( A => operand_a(8), ZN => notA_8_port);
   U74 : INV_X1 port map( A => operand_a(9), ZN => notA_9_port);
   U75 : INV_X1 port map( A => operand_a(10), ZN => notA_10_port);
   U76 : INV_X1 port map( A => operand_a(11), ZN => notA_11_port);
   U77 : INV_X1 port map( A => operand_a(12), ZN => notA_12_port);
   U78 : INV_X1 port map( A => operand_a(13), ZN => notA_13_port);
   U79 : INV_X1 port map( A => operand_a(14), ZN => notA_14_port);
   U80 : INV_X1 port map( A => operand_a(15), ZN => notA_15_port);
   U81 : INV_X1 port map( A => operand_a(16), ZN => notA_16_port);
   U82 : INV_X1 port map( A => operand_a(17), ZN => notA_17_port);
   U83 : INV_X1 port map( A => operand_a(18), ZN => notA_18_port);
   U84 : INV_X1 port map( A => operand_a(19), ZN => notA_19_port);
   U85 : INV_X1 port map( A => operand_a(20), ZN => notA_20_port);
   U86 : INV_X1 port map( A => operand_a(21), ZN => notA_21_port);
   U87 : INV_X1 port map( A => operand_a(22), ZN => notA_22_port);
   U88 : INV_X1 port map( A => operand_a(23), ZN => notA_23_port);
   U89 : INV_X1 port map( A => operand_a(24), ZN => notA_24_port);
   U90 : INV_X1 port map( A => operand_a(25), ZN => notA_25_port);
   U91 : INV_X1 port map( A => operand_a(26), ZN => notA_26_port);
   U92 : INV_X1 port map( A => operand_a(27), ZN => notA_27_port);
   U93 : INV_X1 port map( A => operand_a(28), ZN => notA_28_port);
   U94 : INV_X1 port map( A => operand_a(29), ZN => notA_29_port);
   U95 : INV_X1 port map( A => operand_a(30), ZN => notA_30_port);
   U96 : INV_X1 port map( A => operand_a(31), ZN => notA_31_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity mux5x1 is

   port( a, b, c, d, e : in std_logic_vector (31 downto 0);  enable : in 
         std_logic;  sel : in std_logic_vector (2 downto 0);  out_res : out 
         std_logic_vector (31 downto 0));

end mux5x1;

architecture SYN_Behavioral of mux5x1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n138, n4, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n73, n74, n75, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230 : std_logic;

begin
   
   out_res_tri_8_inst : TBUF_X1 port map( A => n128, EN => n228, Z => 
                           out_res(8));
   out_res_tri_9_inst : TBUF_X1 port map( A => n126, EN => n228, Z => 
                           out_res(9));
   out_res_tri_10_inst : TBUF_X1 port map( A => n125, EN => n228, Z => 
                           out_res(10));
   out_res_tri_11_inst : TBUF_X1 port map( A => n124, EN => n228, Z => 
                           out_res(11));
   out_res_tri_12_inst : TBUF_X1 port map( A => n123, EN => n228, Z => 
                           out_res(12));
   out_res_tri_13_inst : TBUF_X1 port map( A => n122, EN => n228, Z => 
                           out_res(13));
   out_res_tri_14_inst : TBUF_X1 port map( A => n121, EN => n228, Z => 
                           out_res(14));
   out_res_tri_15_inst : TBUF_X1 port map( A => n120, EN => n228, Z => 
                           out_res(15));
   out_res_tri_16_inst : TBUF_X1 port map( A => n119, EN => n226, Z => 
                           out_res(16));
   out_res_tri_17_inst : TBUF_X1 port map( A => n118, EN => n226, Z => 
                           out_res(17));
   out_res_tri_18_inst : TBUF_X1 port map( A => n117, EN => n226, Z => 
                           out_res(18));
   out_res_tri_19_inst : TBUF_X1 port map( A => n116, EN => n226, Z => 
                           out_res(19));
   out_res_tri_20_inst : TBUF_X1 port map( A => n115, EN => n226, Z => 
                           out_res(20));
   out_res_tri_21_inst : TBUF_X1 port map( A => n114, EN => n226, Z => 
                           out_res(21));
   out_res_tri_22_inst : TBUF_X1 port map( A => n113, EN => n226, Z => 
                           out_res(22));
   out_res_tri_23_inst : TBUF_X1 port map( A => n112, EN => n226, Z => 
                           out_res(23));
   out_res_tri_24_inst : TBUF_X1 port map( A => n111, EN => n226, Z => 
                           out_res(24));
   out_res_tri_25_inst : TBUF_X1 port map( A => n110, EN => n226, Z => 
                           out_res(25));
   out_res_tri_26_inst : TBUF_X1 port map( A => n109, EN => n226, Z => 
                           out_res(26));
   out_res_tri_27_inst : TBUF_X1 port map( A => n108, EN => n226, Z => 
                           out_res(27));
   out_res_tri_28_inst : TBUF_X1 port map( A => n107, EN => n227, Z => 
                           out_res(28));
   out_res_tri_29_inst : TBUF_X1 port map( A => n106, EN => n227, Z => 
                           out_res(29));
   out_res_tri_30_inst : TBUF_X1 port map( A => n105, EN => n227, Z => 
                           out_res(30));
   out_res_tri_31_inst : TBUF_X1 port map( A => n104, EN => n227, Z => 
                           out_res(31));
   out_res_tri_0_inst : TBUF_X1 port map( A => n136, EN => n227, Z => 
                           out_res(0));
   out_res_tri_1_inst : TBUF_X1 port map( A => n135, EN => n227, Z => 
                           out_res(1));
   out_res_tri_2_inst : TBUF_X1 port map( A => n134, EN => n227, Z => 
                           out_res(2));
   out_res_tri_3_inst : TBUF_X1 port map( A => n133, EN => n227, Z => 
                           out_res(3));
   out_res_tri_4_inst : TBUF_X1 port map( A => n132, EN => n227, Z => 
                           out_res(4));
   out_res_tri_5_inst : TBUF_X1 port map( A => n131, EN => n227, Z => 
                           out_res(5));
   out_res_tri_6_inst : TBUF_X1 port map( A => n130, EN => n227, Z => 
                           out_res(6));
   out_res_tri_7_inst : TBUF_X1 port map( A => n129, EN => n227, Z => 
                           out_res(7));
   U2 : INV_X1 port map( A => n230, ZN => n229);
   U3 : BUF_X1 port map( A => n11, Z => n214);
   U4 : BUF_X1 port map( A => n11, Z => n215);
   U5 : BUF_X1 port map( A => n10, Z => n217);
   U6 : BUF_X1 port map( A => n10, Z => n218);
   U7 : BUF_X1 port map( A => n8, Z => n223);
   U8 : BUF_X1 port map( A => n8, Z => n224);
   U9 : BUF_X1 port map( A => n10, Z => n219);
   U10 : BUF_X1 port map( A => n11, Z => n216);
   U11 : BUF_X1 port map( A => n8, Z => n225);
   U12 : NOR2_X1 port map( A1 => n74, A2 => sel(0), ZN => n10);
   U13 : BUF_X1 port map( A => n9, Z => n220);
   U14 : BUF_X1 port map( A => n9, Z => n221);
   U15 : NOR2_X1 port map( A1 => n74, A2 => n75, ZN => n8);
   U16 : BUF_X1 port map( A => n9, Z => n222);
   U17 : INV_X1 port map( A => sel(0), ZN => n75);
   U18 : AND2_X1 port map( A1 => n4, A2 => n230, ZN => n11);
   U19 : BUF_X1 port map( A => n138, Z => n227);
   U20 : BUF_X1 port map( A => n138, Z => n226);
   U21 : NOR2_X1 port map( A1 => n75, A2 => sel(1), ZN => n9);
   U22 : NOR2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n4);
   U23 : BUF_X1 port map( A => n138, Z => n228);
   U24 : INV_X1 port map( A => sel(1), ZN => n74);
   U25 : OAI21_X1 port map( B1 => n4, B2 => n230, A => enable, ZN => n138);
   U26 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => n136);
   U27 : AOI222_X1 port map( A1 => d(0), A2 => n225, B1 => b(0), B2 => n222, C1
                           => c(0), C2 => n219, ZN => n7);
   U28 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => n129);
   U29 : AOI22_X1 port map( A1 => a(7), A2 => n216, B1 => e(7), B2 => sel(2), 
                           ZN => n24);
   U30 : AOI222_X1 port map( A1 => d(7), A2 => n225, B1 => b(7), B2 => n222, C1
                           => c(7), C2 => n219, ZN => n25);
   U31 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => n130);
   U32 : AOI22_X1 port map( A1 => a(6), A2 => n216, B1 => e(6), B2 => sel(2), 
                           ZN => n22);
   U33 : AOI222_X1 port map( A1 => d(6), A2 => n225, B1 => b(6), B2 => n222, C1
                           => c(6), C2 => n219, ZN => n23);
   U34 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n131);
   U35 : AOI22_X1 port map( A1 => a(5), A2 => n216, B1 => e(5), B2 => sel(2), 
                           ZN => n20);
   U36 : AOI222_X1 port map( A1 => d(5), A2 => n225, B1 => b(5), B2 => n222, C1
                           => c(5), C2 => n219, ZN => n21);
   U37 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => n132);
   U38 : AOI22_X1 port map( A1 => a(4), A2 => n216, B1 => e(4), B2 => sel(2), 
                           ZN => n18);
   U39 : AOI222_X1 port map( A1 => d(4), A2 => n225, B1 => b(4), B2 => n222, C1
                           => c(4), C2 => n219, ZN => n19);
   U40 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n133);
   U41 : AOI22_X1 port map( A1 => a(3), A2 => n216, B1 => e(3), B2 => sel(2), 
                           ZN => n16);
   U42 : AOI222_X1 port map( A1 => d(3), A2 => n225, B1 => b(3), B2 => n222, C1
                           => c(3), C2 => n219, ZN => n17);
   U43 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n134);
   U44 : AOI22_X1 port map( A1 => a(2), A2 => n216, B1 => e(2), B2 => sel(2), 
                           ZN => n14);
   U45 : AOI222_X1 port map( A1 => d(2), A2 => n225, B1 => b(2), B2 => n222, C1
                           => c(2), C2 => n219, ZN => n15);
   U46 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => n135);
   U47 : AOI22_X1 port map( A1 => a(1), A2 => n216, B1 => e(1), B2 => sel(2), 
                           ZN => n12);
   U48 : AOI222_X1 port map( A1 => d(1), A2 => n225, B1 => b(1), B2 => n222, C1
                           => c(1), C2 => n219, ZN => n13);
   U49 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => n120);
   U50 : AOI22_X1 port map( A1 => a(15), A2 => n215, B1 => e(15), B2 => sel(2),
                           ZN => n40);
   U51 : AOI222_X1 port map( A1 => d(15), A2 => n224, B1 => b(15), B2 => n221, 
                           C1 => c(15), C2 => n218, ZN => n41);
   U52 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => n121);
   U53 : AOI22_X1 port map( A1 => a(14), A2 => n215, B1 => e(14), B2 => n229, 
                           ZN => n38);
   U54 : AOI222_X1 port map( A1 => d(14), A2 => n224, B1 => b(14), B2 => n221, 
                           C1 => c(14), C2 => n218, ZN => n39);
   U55 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => n122);
   U56 : AOI22_X1 port map( A1 => a(13), A2 => n215, B1 => e(13), B2 => sel(2),
                           ZN => n36);
   U57 : AOI222_X1 port map( A1 => d(13), A2 => n224, B1 => b(13), B2 => n221, 
                           C1 => c(13), C2 => n218, ZN => n37);
   U58 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => n123);
   U59 : AOI22_X1 port map( A1 => a(12), A2 => n215, B1 => e(12), B2 => n229, 
                           ZN => n34);
   U60 : AOI222_X1 port map( A1 => d(12), A2 => n224, B1 => b(12), B2 => n221, 
                           C1 => c(12), C2 => n218, ZN => n35);
   U61 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => n124);
   U62 : AOI22_X1 port map( A1 => a(11), A2 => n215, B1 => e(11), B2 => sel(2),
                           ZN => n32);
   U63 : AOI222_X1 port map( A1 => d(11), A2 => n224, B1 => b(11), B2 => n221, 
                           C1 => c(11), C2 => n218, ZN => n33);
   U64 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => n125);
   U65 : AOI22_X1 port map( A1 => a(10), A2 => n215, B1 => e(10), B2 => n229, 
                           ZN => n30);
   U66 : AOI222_X1 port map( A1 => d(10), A2 => n224, B1 => b(10), B2 => n221, 
                           C1 => c(10), C2 => n218, ZN => n31);
   U67 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n126);
   U68 : AOI22_X1 port map( A1 => a(9), A2 => n215, B1 => e(9), B2 => sel(2), 
                           ZN => n28);
   U69 : AOI222_X1 port map( A1 => d(9), A2 => n224, B1 => b(9), B2 => n221, C1
                           => c(9), C2 => n218, ZN => n29);
   U70 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n128);
   U71 : AOI22_X1 port map( A1 => a(8), A2 => n215, B1 => e(8), B2 => n229, ZN 
                           => n26);
   U72 : AOI222_X1 port map( A1 => d(8), A2 => n224, B1 => b(8), B2 => n221, C1
                           => c(8), C2 => n218, ZN => n27);
   U73 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => n104);
   U74 : AOI22_X1 port map( A1 => a(31), A2 => n214, B1 => e(31), B2 => n229, 
                           ZN => n72);
   U75 : AOI222_X1 port map( A1 => d(31), A2 => n223, B1 => b(31), B2 => n220, 
                           C1 => c(31), C2 => n217, ZN => n73);
   U76 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => n105);
   U77 : AOI22_X1 port map( A1 => a(30), A2 => n214, B1 => e(30), B2 => n229, 
                           ZN => n70);
   U78 : AOI222_X1 port map( A1 => d(30), A2 => n223, B1 => b(30), B2 => n220, 
                           C1 => c(30), C2 => n217, ZN => n71);
   U79 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => n106);
   U80 : AOI22_X1 port map( A1 => a(29), A2 => n214, B1 => e(29), B2 => n229, 
                           ZN => n68);
   U81 : AOI222_X1 port map( A1 => d(29), A2 => n223, B1 => b(29), B2 => n220, 
                           C1 => c(29), C2 => n217, ZN => n69);
   U82 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => n107);
   U83 : AOI22_X1 port map( A1 => a(28), A2 => n214, B1 => e(28), B2 => n229, 
                           ZN => n66);
   U84 : AOI222_X1 port map( A1 => d(28), A2 => n223, B1 => b(28), B2 => n220, 
                           C1 => c(28), C2 => n217, ZN => n67);
   U85 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => n108);
   U86 : AOI22_X1 port map( A1 => a(27), A2 => n214, B1 => e(27), B2 => n229, 
                           ZN => n64);
   U87 : AOI222_X1 port map( A1 => d(27), A2 => n223, B1 => b(27), B2 => n220, 
                           C1 => c(27), C2 => n217, ZN => n65);
   U88 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => n109);
   U89 : AOI22_X1 port map( A1 => a(26), A2 => n214, B1 => e(26), B2 => n229, 
                           ZN => n62);
   U90 : AOI222_X1 port map( A1 => d(26), A2 => n223, B1 => b(26), B2 => n220, 
                           C1 => c(26), C2 => n217, ZN => n63);
   U91 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n110);
   U92 : AOI22_X1 port map( A1 => a(25), A2 => n214, B1 => e(25), B2 => n229, 
                           ZN => n60);
   U93 : AOI222_X1 port map( A1 => d(25), A2 => n223, B1 => b(25), B2 => n220, 
                           C1 => c(25), C2 => n217, ZN => n61);
   U94 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => n111);
   U95 : AOI22_X1 port map( A1 => a(24), A2 => n214, B1 => e(24), B2 => n229, 
                           ZN => n58);
   U96 : AOI222_X1 port map( A1 => d(24), A2 => n223, B1 => b(24), B2 => n220, 
                           C1 => c(24), C2 => n217, ZN => n59);
   U97 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => n112);
   U98 : AOI22_X1 port map( A1 => a(23), A2 => n214, B1 => e(23), B2 => n229, 
                           ZN => n56);
   U99 : AOI222_X1 port map( A1 => d(23), A2 => n223, B1 => b(23), B2 => n220, 
                           C1 => c(23), C2 => n217, ZN => n57);
   U100 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => n113);
   U101 : AOI22_X1 port map( A1 => a(22), A2 => n214, B1 => e(22), B2 => n229, 
                           ZN => n54);
   U102 : AOI222_X1 port map( A1 => d(22), A2 => n223, B1 => b(22), B2 => n220,
                           C1 => c(22), C2 => n217, ZN => n55);
   U103 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => n114);
   U104 : AOI22_X1 port map( A1 => a(21), A2 => n214, B1 => e(21), B2 => n229, 
                           ZN => n52);
   U105 : AOI222_X1 port map( A1 => d(21), A2 => n223, B1 => b(21), B2 => n220,
                           C1 => c(21), C2 => n217, ZN => n53);
   U106 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => n115);
   U107 : AOI22_X1 port map( A1 => a(20), A2 => n214, B1 => e(20), B2 => n229, 
                           ZN => n50);
   U108 : AOI222_X1 port map( A1 => d(20), A2 => n223, B1 => b(20), B2 => n220,
                           C1 => c(20), C2 => n217, ZN => n51);
   U109 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => n116);
   U110 : AOI22_X1 port map( A1 => a(19), A2 => n215, B1 => e(19), B2 => sel(2)
                           , ZN => n48);
   U111 : AOI222_X1 port map( A1 => d(19), A2 => n224, B1 => b(19), B2 => n221,
                           C1 => c(19), C2 => n218, ZN => n49);
   U112 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => n117);
   U113 : AOI22_X1 port map( A1 => a(18), A2 => n215, B1 => e(18), B2 => n229, 
                           ZN => n46);
   U114 : AOI222_X1 port map( A1 => d(18), A2 => n224, B1 => b(18), B2 => n221,
                           C1 => c(18), C2 => n218, ZN => n47);
   U115 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n118);
   U116 : AOI22_X1 port map( A1 => a(17), A2 => n215, B1 => e(17), B2 => sel(2)
                           , ZN => n44);
   U117 : AOI222_X1 port map( A1 => d(17), A2 => n224, B1 => b(17), B2 => n221,
                           C1 => c(17), C2 => n218, ZN => n45);
   U118 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => n119);
   U119 : AOI22_X1 port map( A1 => a(16), A2 => n215, B1 => e(16), B2 => n229, 
                           ZN => n42);
   U120 : AOI222_X1 port map( A1 => d(16), A2 => n224, B1 => b(16), B2 => n221,
                           C1 => c(16), C2 => n218, ZN => n43);
   U121 : AOI22_X1 port map( A1 => a(0), A2 => n216, B1 => e(0), B2 => n229, ZN
                           => n6);
   U122 : INV_X1 port map( A => sel(2), ZN => n230);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity booths_mul_N_bit16 is

   port( multiplier, multiplicand : in std_logic_vector (15 downto 0);  product
         : out std_logic_vector (31 downto 0));

end booths_mul_N_bit16;

architecture SYN_Structural of booths_mul_N_bit16 is

   component pentium4_adder_XBIT32_NBIT4_1
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component generator_N_bit16_1
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_2
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component generator_N_bit16_2
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_3
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component generator_N_bit16_3
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_4
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component generator_N_bit16_4
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_5
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component generator_N_bit16_5
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_6
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component generator_N_bit16_6
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_7
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component generator_N_bit16_7
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   component generator_N_bit16_0
      port( multiplicant : in std_logic_vector (15 downto 0);  N_shift : in 
            std_logic_vector (0 to 31);  select_signal : in std_logic_vector (2
            downto 0);  Out_value : out std_logic_vector (31 downto 0));
   end component;
   
   signal routing_wires_9_9_port, routing_wires_9_8_port, 
      routing_wires_9_7_port, routing_wires_9_6_port, routing_wires_9_5_port, 
      routing_wires_9_4_port, routing_wires_9_3_port, routing_wires_9_31_port, 
      routing_wires_9_30_port, routing_wires_9_2_port, routing_wires_9_29_port,
      routing_wires_9_28_port, routing_wires_9_27_port, routing_wires_9_26_port
      , routing_wires_9_25_port, routing_wires_9_24_port, 
      routing_wires_9_23_port, routing_wires_9_22_port, routing_wires_9_21_port
      , routing_wires_9_20_port, routing_wires_9_1_port, 
      routing_wires_9_19_port, routing_wires_9_18_port, routing_wires_9_17_port
      , routing_wires_9_16_port, routing_wires_9_15_port, 
      routing_wires_9_14_port, routing_wires_9_13_port, routing_wires_9_12_port
      , routing_wires_9_11_port, routing_wires_9_10_port, 
      routing_wires_9_0_port, routing_wires_8_9_port, routing_wires_8_8_port, 
      routing_wires_8_7_port, routing_wires_8_6_port, routing_wires_8_5_port, 
      routing_wires_8_4_port, routing_wires_8_3_port, routing_wires_8_31_port, 
      routing_wires_8_30_port, routing_wires_8_2_port, routing_wires_8_29_port,
      routing_wires_8_28_port, routing_wires_8_27_port, routing_wires_8_26_port
      , routing_wires_8_25_port, routing_wires_8_24_port, 
      routing_wires_8_23_port, routing_wires_8_22_port, routing_wires_8_21_port
      , routing_wires_8_20_port, routing_wires_8_1_port, 
      routing_wires_8_19_port, routing_wires_8_18_port, routing_wires_8_17_port
      , routing_wires_8_16_port, routing_wires_8_15_port, 
      routing_wires_8_14_port, routing_wires_8_13_port, routing_wires_8_12_port
      , routing_wires_8_11_port, routing_wires_8_10_port, 
      routing_wires_8_0_port, routing_wires_7_9_port, routing_wires_7_8_port, 
      routing_wires_7_7_port, routing_wires_7_6_port, routing_wires_7_5_port, 
      routing_wires_7_4_port, routing_wires_7_3_port, routing_wires_7_31_port, 
      routing_wires_7_30_port, routing_wires_7_2_port, routing_wires_7_29_port,
      routing_wires_7_28_port, routing_wires_7_27_port, routing_wires_7_26_port
      , routing_wires_7_25_port, routing_wires_7_24_port, 
      routing_wires_7_23_port, routing_wires_7_22_port, routing_wires_7_21_port
      , routing_wires_7_20_port, routing_wires_7_1_port, 
      routing_wires_7_19_port, routing_wires_7_18_port, routing_wires_7_17_port
      , routing_wires_7_16_port, routing_wires_7_15_port, 
      routing_wires_7_14_port, routing_wires_7_13_port, routing_wires_7_12_port
      , routing_wires_7_11_port, routing_wires_7_10_port, 
      routing_wires_7_0_port, routing_wires_6_9_port, routing_wires_6_8_port, 
      routing_wires_6_7_port, routing_wires_6_6_port, routing_wires_6_5_port, 
      routing_wires_6_4_port, routing_wires_6_3_port, routing_wires_6_31_port, 
      routing_wires_6_30_port, routing_wires_6_2_port, routing_wires_6_29_port,
      routing_wires_6_28_port, routing_wires_6_27_port, routing_wires_6_26_port
      , routing_wires_6_25_port, routing_wires_6_24_port, 
      routing_wires_6_23_port, routing_wires_6_22_port, routing_wires_6_21_port
      , routing_wires_6_20_port, routing_wires_6_1_port, 
      routing_wires_6_19_port, routing_wires_6_18_port, routing_wires_6_17_port
      , routing_wires_6_16_port, routing_wires_6_15_port, 
      routing_wires_6_14_port, routing_wires_6_13_port, routing_wires_6_12_port
      , routing_wires_6_11_port, routing_wires_6_10_port, 
      routing_wires_6_0_port, routing_wires_5_9_port, routing_wires_5_8_port, 
      routing_wires_5_7_port, routing_wires_5_6_port, routing_wires_5_5_port, 
      routing_wires_5_4_port, routing_wires_5_3_port, routing_wires_5_31_port, 
      routing_wires_5_30_port, routing_wires_5_2_port, routing_wires_5_29_port,
      routing_wires_5_28_port, routing_wires_5_27_port, routing_wires_5_26_port
      , routing_wires_5_25_port, routing_wires_5_24_port, 
      routing_wires_5_23_port, routing_wires_5_22_port, routing_wires_5_21_port
      , routing_wires_5_20_port, routing_wires_5_1_port, 
      routing_wires_5_19_port, routing_wires_5_18_port, routing_wires_5_17_port
      , routing_wires_5_16_port, routing_wires_5_15_port, 
      routing_wires_5_14_port, routing_wires_5_13_port, routing_wires_5_12_port
      , routing_wires_5_11_port, routing_wires_5_10_port, 
      routing_wires_5_0_port, routing_wires_4_9_port, routing_wires_4_8_port, 
      routing_wires_4_7_port, routing_wires_4_6_port, routing_wires_4_5_port, 
      routing_wires_4_4_port, routing_wires_4_3_port, routing_wires_4_31_port, 
      routing_wires_4_30_port, routing_wires_4_2_port, routing_wires_4_29_port,
      routing_wires_4_28_port, routing_wires_4_27_port, routing_wires_4_26_port
      , routing_wires_4_25_port, routing_wires_4_24_port, 
      routing_wires_4_23_port, routing_wires_4_22_port, routing_wires_4_21_port
      , routing_wires_4_20_port, routing_wires_4_1_port, 
      routing_wires_4_19_port, routing_wires_4_18_port, routing_wires_4_17_port
      , routing_wires_4_16_port, routing_wires_4_15_port, 
      routing_wires_4_14_port, routing_wires_4_13_port, routing_wires_4_12_port
      , routing_wires_4_11_port, routing_wires_4_10_port, 
      routing_wires_4_0_port, routing_wires_3_9_port, routing_wires_3_8_port, 
      routing_wires_3_7_port, routing_wires_3_6_port, routing_wires_3_5_port, 
      routing_wires_3_4_port, routing_wires_3_3_port, routing_wires_3_31_port, 
      routing_wires_3_30_port, routing_wires_3_2_port, routing_wires_3_29_port,
      routing_wires_3_28_port, routing_wires_3_27_port, routing_wires_3_26_port
      , routing_wires_3_25_port, routing_wires_3_24_port, 
      routing_wires_3_23_port, routing_wires_3_22_port, routing_wires_3_21_port
      , routing_wires_3_20_port, routing_wires_3_1_port, 
      routing_wires_3_19_port, routing_wires_3_18_port, routing_wires_3_17_port
      , routing_wires_3_16_port, routing_wires_3_15_port, 
      routing_wires_3_14_port, routing_wires_3_13_port, routing_wires_3_12_port
      , routing_wires_3_11_port, routing_wires_3_10_port, 
      routing_wires_3_0_port, routing_wires_2_9_port, routing_wires_2_8_port, 
      routing_wires_2_7_port, routing_wires_2_6_port, routing_wires_2_5_port, 
      routing_wires_2_4_port, routing_wires_2_3_port, routing_wires_2_31_port, 
      routing_wires_2_30_port, routing_wires_2_2_port, routing_wires_2_29_port,
      routing_wires_2_28_port, routing_wires_2_27_port, routing_wires_2_26_port
      , routing_wires_2_25_port, routing_wires_2_24_port, 
      routing_wires_2_23_port, routing_wires_2_22_port, routing_wires_2_21_port
      , routing_wires_2_20_port, routing_wires_2_1_port, 
      routing_wires_2_19_port, routing_wires_2_18_port, routing_wires_2_17_port
      , routing_wires_2_16_port, routing_wires_2_15_port, 
      routing_wires_2_14_port, routing_wires_2_13_port, routing_wires_2_12_port
      , routing_wires_2_11_port, routing_wires_2_10_port, 
      routing_wires_2_0_port, routing_wires_1_9_port, routing_wires_1_8_port, 
      routing_wires_1_7_port, routing_wires_1_6_port, routing_wires_1_5_port, 
      routing_wires_1_4_port, routing_wires_1_3_port, routing_wires_1_31_port, 
      routing_wires_1_30_port, routing_wires_1_2_port, routing_wires_1_29_port,
      routing_wires_1_28_port, routing_wires_1_27_port, routing_wires_1_26_port
      , routing_wires_1_25_port, routing_wires_1_24_port, 
      routing_wires_1_23_port, routing_wires_1_22_port, routing_wires_1_21_port
      , routing_wires_1_20_port, routing_wires_1_1_port, 
      routing_wires_1_19_port, routing_wires_1_18_port, routing_wires_1_17_port
      , routing_wires_1_16_port, routing_wires_1_15_port, 
      routing_wires_1_14_port, routing_wires_1_13_port, routing_wires_1_12_port
      , routing_wires_1_11_port, routing_wires_1_10_port, 
      routing_wires_1_0_port, routing_wires_14_9_port, routing_wires_14_8_port,
      routing_wires_14_7_port, routing_wires_14_6_port, routing_wires_14_5_port
      , routing_wires_14_4_port, routing_wires_14_3_port, 
      routing_wires_14_31_port, routing_wires_14_30_port, 
      routing_wires_14_2_port, routing_wires_14_29_port, 
      routing_wires_14_28_port, routing_wires_14_27_port, 
      routing_wires_14_26_port, routing_wires_14_25_port, 
      routing_wires_14_24_port, routing_wires_14_23_port, 
      routing_wires_14_22_port, routing_wires_14_21_port, 
      routing_wires_14_20_port, routing_wires_14_1_port, 
      routing_wires_14_19_port, routing_wires_14_18_port, 
      routing_wires_14_17_port, routing_wires_14_16_port, 
      routing_wires_14_15_port, routing_wires_14_14_port, 
      routing_wires_14_13_port, routing_wires_14_12_port, 
      routing_wires_14_11_port, routing_wires_14_10_port, 
      routing_wires_14_0_port, routing_wires_13_9_port, routing_wires_13_8_port
      , routing_wires_13_7_port, routing_wires_13_6_port, 
      routing_wires_13_5_port, routing_wires_13_4_port, routing_wires_13_3_port
      , routing_wires_13_31_port, routing_wires_13_30_port, 
      routing_wires_13_2_port, routing_wires_13_29_port, 
      routing_wires_13_28_port, routing_wires_13_27_port, 
      routing_wires_13_26_port, routing_wires_13_25_port, 
      routing_wires_13_24_port, routing_wires_13_23_port, 
      routing_wires_13_22_port, routing_wires_13_21_port, 
      routing_wires_13_20_port, routing_wires_13_1_port, 
      routing_wires_13_19_port, routing_wires_13_18_port, 
      routing_wires_13_17_port, routing_wires_13_16_port, 
      routing_wires_13_15_port, routing_wires_13_14_port, 
      routing_wires_13_13_port, routing_wires_13_12_port, 
      routing_wires_13_11_port, routing_wires_13_10_port, 
      routing_wires_13_0_port, routing_wires_12_9_port, routing_wires_12_8_port
      , routing_wires_12_7_port, routing_wires_12_6_port, 
      routing_wires_12_5_port, routing_wires_12_4_port, routing_wires_12_3_port
      , routing_wires_12_31_port, routing_wires_12_30_port, 
      routing_wires_12_2_port, routing_wires_12_29_port, 
      routing_wires_12_28_port, routing_wires_12_27_port, 
      routing_wires_12_26_port, routing_wires_12_25_port, 
      routing_wires_12_24_port, routing_wires_12_23_port, 
      routing_wires_12_22_port, routing_wires_12_21_port, 
      routing_wires_12_20_port, routing_wires_12_1_port, 
      routing_wires_12_19_port, routing_wires_12_18_port, 
      routing_wires_12_17_port, routing_wires_12_16_port, 
      routing_wires_12_15_port, routing_wires_12_14_port, 
      routing_wires_12_13_port, routing_wires_12_12_port, 
      routing_wires_12_11_port, routing_wires_12_10_port, 
      routing_wires_12_0_port, routing_wires_11_9_port, routing_wires_11_8_port
      , routing_wires_11_7_port, routing_wires_11_6_port, 
      routing_wires_11_5_port, routing_wires_11_4_port, routing_wires_11_3_port
      , routing_wires_11_31_port, routing_wires_11_30_port, 
      routing_wires_11_2_port, routing_wires_11_29_port, 
      routing_wires_11_28_port, routing_wires_11_27_port, 
      routing_wires_11_26_port, routing_wires_11_25_port, 
      routing_wires_11_24_port, routing_wires_11_23_port, 
      routing_wires_11_22_port, routing_wires_11_21_port, 
      routing_wires_11_20_port, routing_wires_11_1_port, 
      routing_wires_11_19_port, routing_wires_11_18_port, 
      routing_wires_11_17_port, routing_wires_11_16_port, 
      routing_wires_11_15_port, routing_wires_11_14_port, 
      routing_wires_11_13_port, routing_wires_11_12_port, 
      routing_wires_11_11_port, routing_wires_11_10_port, 
      routing_wires_11_0_port, routing_wires_10_9_port, routing_wires_10_8_port
      , routing_wires_10_7_port, routing_wires_10_6_port, 
      routing_wires_10_5_port, routing_wires_10_4_port, routing_wires_10_3_port
      , routing_wires_10_31_port, routing_wires_10_30_port, 
      routing_wires_10_2_port, routing_wires_10_29_port, 
      routing_wires_10_28_port, routing_wires_10_27_port, 
      routing_wires_10_26_port, routing_wires_10_25_port, 
      routing_wires_10_24_port, routing_wires_10_23_port, 
      routing_wires_10_22_port, routing_wires_10_21_port, 
      routing_wires_10_20_port, routing_wires_10_1_port, 
      routing_wires_10_19_port, routing_wires_10_18_port, 
      routing_wires_10_17_port, routing_wires_10_16_port, 
      routing_wires_10_15_port, routing_wires_10_14_port, 
      routing_wires_10_13_port, routing_wires_10_12_port, 
      routing_wires_10_11_port, routing_wires_10_10_port, 
      routing_wires_10_0_port, net3150, net3149, net3148, net3147, net3146, 
      net3145, net3144, n21, n22 : std_logic;
   
   signal N_shift_pin, N_shift_pin_port, N_shift_pin_port2, N_shift_pin_port3, 
      N_shift_pin_port4, N_shift_pin_port5, N_shift_pin_port6, 
      N_shift_pin_port7 : std_logic_vector (0 to 31);

begin
   
   N_shift_pin <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21,
      n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n21 );
   g0_0 : generator_N_bit16_0 port map( multiplicant(15) => multiplicand(15), 
      multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin, select_signal(2) => multiplier(1), 
      select_signal(1) => multiplier(0), select_signal(0) => n21, Out_value(31)
      => routing_wires_1_31_port, Out_value(30) => routing_wires_1_30_port, 
      Out_value(29) => routing_wires_1_29_port, Out_value(28) => 
      routing_wires_1_28_port, Out_value(27) => routing_wires_1_27_port, 
      Out_value(26) => routing_wires_1_26_port, Out_value(25) => 
      routing_wires_1_25_port, Out_value(24) => routing_wires_1_24_port, 
      Out_value(23) => routing_wires_1_23_port, Out_value(22) => 
      routing_wires_1_22_port, Out_value(21) => routing_wires_1_21_port, 
      Out_value(20) => routing_wires_1_20_port, Out_value(19) => 
      routing_wires_1_19_port, Out_value(18) => routing_wires_1_18_port, 
      Out_value(17) => routing_wires_1_17_port, Out_value(16) => 
      routing_wires_1_16_port, Out_value(15) => routing_wires_1_15_port, 
      Out_value(14) => routing_wires_1_14_port, Out_value(13) => 
      routing_wires_1_13_port, Out_value(12) => routing_wires_1_12_port, 
      Out_value(11) => routing_wires_1_11_port, Out_value(10) => 
      routing_wires_1_10_port, Out_value(9) => routing_wires_1_9_port, 
      Out_value(8) => routing_wires_1_8_port, Out_value(7) => 
      routing_wires_1_7_port, Out_value(6) => routing_wires_1_6_port, 
      Out_value(5) => routing_wires_1_5_port, Out_value(4) => 
      routing_wires_1_4_port, Out_value(3) => routing_wires_1_3_port, 
      Out_value(2) => routing_wires_1_2_port, Out_value(1) => 
      routing_wires_1_1_port, Out_value(0) => routing_wires_1_0_port);
   N_shift_pin_port <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21,
      n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n22, n21 );
   g1_0 : generator_N_bit16_7 port map( multiplicant(15) => multiplicand(15), 
      multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin_port, select_signal(2) => multiplier(3), 
      select_signal(1) => multiplier(2), select_signal(0) => multiplier(1), 
      Out_value(31) => routing_wires_2_31_port, Out_value(30) => 
      routing_wires_2_30_port, Out_value(29) => routing_wires_2_29_port, 
      Out_value(28) => routing_wires_2_28_port, Out_value(27) => 
      routing_wires_2_27_port, Out_value(26) => routing_wires_2_26_port, 
      Out_value(25) => routing_wires_2_25_port, Out_value(24) => 
      routing_wires_2_24_port, Out_value(23) => routing_wires_2_23_port, 
      Out_value(22) => routing_wires_2_22_port, Out_value(21) => 
      routing_wires_2_21_port, Out_value(20) => routing_wires_2_20_port, 
      Out_value(19) => routing_wires_2_19_port, Out_value(18) => 
      routing_wires_2_18_port, Out_value(17) => routing_wires_2_17_port, 
      Out_value(16) => routing_wires_2_16_port, Out_value(15) => 
      routing_wires_2_15_port, Out_value(14) => routing_wires_2_14_port, 
      Out_value(13) => routing_wires_2_13_port, Out_value(12) => 
      routing_wires_2_12_port, Out_value(11) => routing_wires_2_11_port, 
      Out_value(10) => routing_wires_2_10_port, Out_value(9) => 
      routing_wires_2_9_port, Out_value(8) => routing_wires_2_8_port, 
      Out_value(7) => routing_wires_2_7_port, Out_value(6) => 
      routing_wires_2_6_port, Out_value(5) => routing_wires_2_5_port, 
      Out_value(4) => routing_wires_2_4_port, Out_value(3) => 
      routing_wires_2_3_port, Out_value(2) => routing_wires_2_2_port, 
      Out_value(1) => routing_wires_2_1_port, Out_value(0) => 
      routing_wires_2_0_port);
   a0_0 : pentium4_adder_XBIT32_NBIT4_7 port map( A(31) => 
                           routing_wires_1_31_port, A(30) => 
                           routing_wires_1_30_port, A(29) => 
                           routing_wires_1_29_port, A(28) => 
                           routing_wires_1_28_port, A(27) => 
                           routing_wires_1_27_port, A(26) => 
                           routing_wires_1_26_port, A(25) => 
                           routing_wires_1_25_port, A(24) => 
                           routing_wires_1_24_port, A(23) => 
                           routing_wires_1_23_port, A(22) => 
                           routing_wires_1_22_port, A(21) => 
                           routing_wires_1_21_port, A(20) => 
                           routing_wires_1_20_port, A(19) => 
                           routing_wires_1_19_port, A(18) => 
                           routing_wires_1_18_port, A(17) => 
                           routing_wires_1_17_port, A(16) => 
                           routing_wires_1_16_port, A(15) => 
                           routing_wires_1_15_port, A(14) => 
                           routing_wires_1_14_port, A(13) => 
                           routing_wires_1_13_port, A(12) => 
                           routing_wires_1_12_port, A(11) => 
                           routing_wires_1_11_port, A(10) => 
                           routing_wires_1_10_port, A(9) => 
                           routing_wires_1_9_port, A(8) => 
                           routing_wires_1_8_port, A(7) => 
                           routing_wires_1_7_port, A(6) => 
                           routing_wires_1_6_port, A(5) => 
                           routing_wires_1_5_port, A(4) => 
                           routing_wires_1_4_port, A(3) => 
                           routing_wires_1_3_port, A(2) => 
                           routing_wires_1_2_port, A(1) => 
                           routing_wires_1_1_port, A(0) => 
                           routing_wires_1_0_port, B(31) => 
                           routing_wires_2_31_port, B(30) => 
                           routing_wires_2_30_port, B(29) => 
                           routing_wires_2_29_port, B(28) => 
                           routing_wires_2_28_port, B(27) => 
                           routing_wires_2_27_port, B(26) => 
                           routing_wires_2_26_port, B(25) => 
                           routing_wires_2_25_port, B(24) => 
                           routing_wires_2_24_port, B(23) => 
                           routing_wires_2_23_port, B(22) => 
                           routing_wires_2_22_port, B(21) => 
                           routing_wires_2_21_port, B(20) => 
                           routing_wires_2_20_port, B(19) => 
                           routing_wires_2_19_port, B(18) => 
                           routing_wires_2_18_port, B(17) => 
                           routing_wires_2_17_port, B(16) => 
                           routing_wires_2_16_port, B(15) => 
                           routing_wires_2_15_port, B(14) => 
                           routing_wires_2_14_port, B(13) => 
                           routing_wires_2_13_port, B(12) => 
                           routing_wires_2_12_port, B(11) => 
                           routing_wires_2_11_port, B(10) => 
                           routing_wires_2_10_port, B(9) => 
                           routing_wires_2_9_port, B(8) => 
                           routing_wires_2_8_port, B(7) => 
                           routing_wires_2_7_port, B(6) => 
                           routing_wires_2_6_port, B(5) => 
                           routing_wires_2_5_port, B(4) => 
                           routing_wires_2_4_port, B(3) => 
                           routing_wires_2_3_port, B(2) => 
                           routing_wires_2_2_port, B(1) => 
                           routing_wires_2_1_port, B(0) => 
                           routing_wires_2_0_port, C_0 => n21, S(31) => 
                           routing_wires_3_31_port, S(30) => 
                           routing_wires_3_30_port, S(29) => 
                           routing_wires_3_29_port, S(28) => 
                           routing_wires_3_28_port, S(27) => 
                           routing_wires_3_27_port, S(26) => 
                           routing_wires_3_26_port, S(25) => 
                           routing_wires_3_25_port, S(24) => 
                           routing_wires_3_24_port, S(23) => 
                           routing_wires_3_23_port, S(22) => 
                           routing_wires_3_22_port, S(21) => 
                           routing_wires_3_21_port, S(20) => 
                           routing_wires_3_20_port, S(19) => 
                           routing_wires_3_19_port, S(18) => 
                           routing_wires_3_18_port, S(17) => 
                           routing_wires_3_17_port, S(16) => 
                           routing_wires_3_16_port, S(15) => 
                           routing_wires_3_15_port, S(14) => 
                           routing_wires_3_14_port, S(13) => 
                           routing_wires_3_13_port, S(12) => 
                           routing_wires_3_12_port, S(11) => 
                           routing_wires_3_11_port, S(10) => 
                           routing_wires_3_10_port, S(9) => 
                           routing_wires_3_9_port, S(8) => 
                           routing_wires_3_8_port, S(7) => 
                           routing_wires_3_7_port, S(6) => 
                           routing_wires_3_6_port, S(5) => 
                           routing_wires_3_5_port, S(4) => 
                           routing_wires_3_4_port, S(3) => 
                           routing_wires_3_3_port, S(2) => 
                           routing_wires_3_2_port, S(1) => 
                           routing_wires_3_1_port, S(0) => 
                           routing_wires_3_0_port, Cout => net3150);
   N_shift_pin_port2 <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, 
      n21, n21, n21, n21, n22, n21, n21 );
   gi_4 : generator_N_bit16_6 port map( multiplicant(15) => multiplicand(15), 
      multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin_port2, select_signal(2) => multiplier(5), 
      select_signal(1) => multiplier(4), select_signal(0) => multiplier(3), 
      Out_value(31) => routing_wires_4_31_port, Out_value(30) => 
      routing_wires_4_30_port, Out_value(29) => routing_wires_4_29_port, 
      Out_value(28) => routing_wires_4_28_port, Out_value(27) => 
      routing_wires_4_27_port, Out_value(26) => routing_wires_4_26_port, 
      Out_value(25) => routing_wires_4_25_port, Out_value(24) => 
      routing_wires_4_24_port, Out_value(23) => routing_wires_4_23_port, 
      Out_value(22) => routing_wires_4_22_port, Out_value(21) => 
      routing_wires_4_21_port, Out_value(20) => routing_wires_4_20_port, 
      Out_value(19) => routing_wires_4_19_port, Out_value(18) => 
      routing_wires_4_18_port, Out_value(17) => routing_wires_4_17_port, 
      Out_value(16) => routing_wires_4_16_port, Out_value(15) => 
      routing_wires_4_15_port, Out_value(14) => routing_wires_4_14_port, 
      Out_value(13) => routing_wires_4_13_port, Out_value(12) => 
      routing_wires_4_12_port, Out_value(11) => routing_wires_4_11_port, 
      Out_value(10) => routing_wires_4_10_port, Out_value(9) => 
      routing_wires_4_9_port, Out_value(8) => routing_wires_4_8_port, 
      Out_value(7) => routing_wires_4_7_port, Out_value(6) => 
      routing_wires_4_6_port, Out_value(5) => routing_wires_4_5_port, 
      Out_value(4) => routing_wires_4_4_port, Out_value(3) => 
      routing_wires_4_3_port, Out_value(2) => routing_wires_4_2_port, 
      Out_value(1) => routing_wires_4_1_port, Out_value(0) => 
      routing_wires_4_0_port);
   ai_4 : pentium4_adder_XBIT32_NBIT4_6 port map( A(31) => 
                           routing_wires_3_31_port, A(30) => 
                           routing_wires_3_30_port, A(29) => 
                           routing_wires_3_29_port, A(28) => 
                           routing_wires_3_28_port, A(27) => 
                           routing_wires_3_27_port, A(26) => 
                           routing_wires_3_26_port, A(25) => 
                           routing_wires_3_25_port, A(24) => 
                           routing_wires_3_24_port, A(23) => 
                           routing_wires_3_23_port, A(22) => 
                           routing_wires_3_22_port, A(21) => 
                           routing_wires_3_21_port, A(20) => 
                           routing_wires_3_20_port, A(19) => 
                           routing_wires_3_19_port, A(18) => 
                           routing_wires_3_18_port, A(17) => 
                           routing_wires_3_17_port, A(16) => 
                           routing_wires_3_16_port, A(15) => 
                           routing_wires_3_15_port, A(14) => 
                           routing_wires_3_14_port, A(13) => 
                           routing_wires_3_13_port, A(12) => 
                           routing_wires_3_12_port, A(11) => 
                           routing_wires_3_11_port, A(10) => 
                           routing_wires_3_10_port, A(9) => 
                           routing_wires_3_9_port, A(8) => 
                           routing_wires_3_8_port, A(7) => 
                           routing_wires_3_7_port, A(6) => 
                           routing_wires_3_6_port, A(5) => 
                           routing_wires_3_5_port, A(4) => 
                           routing_wires_3_4_port, A(3) => 
                           routing_wires_3_3_port, A(2) => 
                           routing_wires_3_2_port, A(1) => 
                           routing_wires_3_1_port, A(0) => 
                           routing_wires_3_0_port, B(31) => 
                           routing_wires_4_31_port, B(30) => 
                           routing_wires_4_30_port, B(29) => 
                           routing_wires_4_29_port, B(28) => 
                           routing_wires_4_28_port, B(27) => 
                           routing_wires_4_27_port, B(26) => 
                           routing_wires_4_26_port, B(25) => 
                           routing_wires_4_25_port, B(24) => 
                           routing_wires_4_24_port, B(23) => 
                           routing_wires_4_23_port, B(22) => 
                           routing_wires_4_22_port, B(21) => 
                           routing_wires_4_21_port, B(20) => 
                           routing_wires_4_20_port, B(19) => 
                           routing_wires_4_19_port, B(18) => 
                           routing_wires_4_18_port, B(17) => 
                           routing_wires_4_17_port, B(16) => 
                           routing_wires_4_16_port, B(15) => 
                           routing_wires_4_15_port, B(14) => 
                           routing_wires_4_14_port, B(13) => 
                           routing_wires_4_13_port, B(12) => 
                           routing_wires_4_12_port, B(11) => 
                           routing_wires_4_11_port, B(10) => 
                           routing_wires_4_10_port, B(9) => 
                           routing_wires_4_9_port, B(8) => 
                           routing_wires_4_8_port, B(7) => 
                           routing_wires_4_7_port, B(6) => 
                           routing_wires_4_6_port, B(5) => 
                           routing_wires_4_5_port, B(4) => 
                           routing_wires_4_4_port, B(3) => 
                           routing_wires_4_3_port, B(2) => 
                           routing_wires_4_2_port, B(1) => 
                           routing_wires_4_1_port, B(0) => 
                           routing_wires_4_0_port, C_0 => n21, S(31) => 
                           routing_wires_5_31_port, S(30) => 
                           routing_wires_5_30_port, S(29) => 
                           routing_wires_5_29_port, S(28) => 
                           routing_wires_5_28_port, S(27) => 
                           routing_wires_5_27_port, S(26) => 
                           routing_wires_5_26_port, S(25) => 
                           routing_wires_5_25_port, S(24) => 
                           routing_wires_5_24_port, S(23) => 
                           routing_wires_5_23_port, S(22) => 
                           routing_wires_5_22_port, S(21) => 
                           routing_wires_5_21_port, S(20) => 
                           routing_wires_5_20_port, S(19) => 
                           routing_wires_5_19_port, S(18) => 
                           routing_wires_5_18_port, S(17) => 
                           routing_wires_5_17_port, S(16) => 
                           routing_wires_5_16_port, S(15) => 
                           routing_wires_5_15_port, S(14) => 
                           routing_wires_5_14_port, S(13) => 
                           routing_wires_5_13_port, S(12) => 
                           routing_wires_5_12_port, S(11) => 
                           routing_wires_5_11_port, S(10) => 
                           routing_wires_5_10_port, S(9) => 
                           routing_wires_5_9_port, S(8) => 
                           routing_wires_5_8_port, S(7) => 
                           routing_wires_5_7_port, S(6) => 
                           routing_wires_5_6_port, S(5) => 
                           routing_wires_5_5_port, S(4) => 
                           routing_wires_5_4_port, S(3) => 
                           routing_wires_5_3_port, S(2) => 
                           routing_wires_5_2_port, S(1) => 
                           routing_wires_5_1_port, S(0) => 
                           routing_wires_5_0_port, Cout => net3149);
   N_shift_pin_port3 <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, 
      n21, n21, n21, n21, n22, n22, n21 );
   gi_6 : generator_N_bit16_5 port map( multiplicant(15) => multiplicand(15), 
      multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin_port3, select_signal(2) => multiplier(7), 
      select_signal(1) => multiplier(6), select_signal(0) => multiplier(5), 
      Out_value(31) => routing_wires_6_31_port, Out_value(30) => 
      routing_wires_6_30_port, Out_value(29) => routing_wires_6_29_port, 
      Out_value(28) => routing_wires_6_28_port, Out_value(27) => 
      routing_wires_6_27_port, Out_value(26) => routing_wires_6_26_port, 
      Out_value(25) => routing_wires_6_25_port, Out_value(24) => 
      routing_wires_6_24_port, Out_value(23) => routing_wires_6_23_port, 
      Out_value(22) => routing_wires_6_22_port, Out_value(21) => 
      routing_wires_6_21_port, Out_value(20) => routing_wires_6_20_port, 
      Out_value(19) => routing_wires_6_19_port, Out_value(18) => 
      routing_wires_6_18_port, Out_value(17) => routing_wires_6_17_port, 
      Out_value(16) => routing_wires_6_16_port, Out_value(15) => 
      routing_wires_6_15_port, Out_value(14) => routing_wires_6_14_port, 
      Out_value(13) => routing_wires_6_13_port, Out_value(12) => 
      routing_wires_6_12_port, Out_value(11) => routing_wires_6_11_port, 
      Out_value(10) => routing_wires_6_10_port, Out_value(9) => 
      routing_wires_6_9_port, Out_value(8) => routing_wires_6_8_port, 
      Out_value(7) => routing_wires_6_7_port, Out_value(6) => 
      routing_wires_6_6_port, Out_value(5) => routing_wires_6_5_port, 
      Out_value(4) => routing_wires_6_4_port, Out_value(3) => 
      routing_wires_6_3_port, Out_value(2) => routing_wires_6_2_port, 
      Out_value(1) => routing_wires_6_1_port, Out_value(0) => 
      routing_wires_6_0_port);
   ai_6 : pentium4_adder_XBIT32_NBIT4_5 port map( A(31) => 
                           routing_wires_5_31_port, A(30) => 
                           routing_wires_5_30_port, A(29) => 
                           routing_wires_5_29_port, A(28) => 
                           routing_wires_5_28_port, A(27) => 
                           routing_wires_5_27_port, A(26) => 
                           routing_wires_5_26_port, A(25) => 
                           routing_wires_5_25_port, A(24) => 
                           routing_wires_5_24_port, A(23) => 
                           routing_wires_5_23_port, A(22) => 
                           routing_wires_5_22_port, A(21) => 
                           routing_wires_5_21_port, A(20) => 
                           routing_wires_5_20_port, A(19) => 
                           routing_wires_5_19_port, A(18) => 
                           routing_wires_5_18_port, A(17) => 
                           routing_wires_5_17_port, A(16) => 
                           routing_wires_5_16_port, A(15) => 
                           routing_wires_5_15_port, A(14) => 
                           routing_wires_5_14_port, A(13) => 
                           routing_wires_5_13_port, A(12) => 
                           routing_wires_5_12_port, A(11) => 
                           routing_wires_5_11_port, A(10) => 
                           routing_wires_5_10_port, A(9) => 
                           routing_wires_5_9_port, A(8) => 
                           routing_wires_5_8_port, A(7) => 
                           routing_wires_5_7_port, A(6) => 
                           routing_wires_5_6_port, A(5) => 
                           routing_wires_5_5_port, A(4) => 
                           routing_wires_5_4_port, A(3) => 
                           routing_wires_5_3_port, A(2) => 
                           routing_wires_5_2_port, A(1) => 
                           routing_wires_5_1_port, A(0) => 
                           routing_wires_5_0_port, B(31) => 
                           routing_wires_6_31_port, B(30) => 
                           routing_wires_6_30_port, B(29) => 
                           routing_wires_6_29_port, B(28) => 
                           routing_wires_6_28_port, B(27) => 
                           routing_wires_6_27_port, B(26) => 
                           routing_wires_6_26_port, B(25) => 
                           routing_wires_6_25_port, B(24) => 
                           routing_wires_6_24_port, B(23) => 
                           routing_wires_6_23_port, B(22) => 
                           routing_wires_6_22_port, B(21) => 
                           routing_wires_6_21_port, B(20) => 
                           routing_wires_6_20_port, B(19) => 
                           routing_wires_6_19_port, B(18) => 
                           routing_wires_6_18_port, B(17) => 
                           routing_wires_6_17_port, B(16) => 
                           routing_wires_6_16_port, B(15) => 
                           routing_wires_6_15_port, B(14) => 
                           routing_wires_6_14_port, B(13) => 
                           routing_wires_6_13_port, B(12) => 
                           routing_wires_6_12_port, B(11) => 
                           routing_wires_6_11_port, B(10) => 
                           routing_wires_6_10_port, B(9) => 
                           routing_wires_6_9_port, B(8) => 
                           routing_wires_6_8_port, B(7) => 
                           routing_wires_6_7_port, B(6) => 
                           routing_wires_6_6_port, B(5) => 
                           routing_wires_6_5_port, B(4) => 
                           routing_wires_6_4_port, B(3) => 
                           routing_wires_6_3_port, B(2) => 
                           routing_wires_6_2_port, B(1) => 
                           routing_wires_6_1_port, B(0) => 
                           routing_wires_6_0_port, C_0 => n21, S(31) => 
                           routing_wires_7_31_port, S(30) => 
                           routing_wires_7_30_port, S(29) => 
                           routing_wires_7_29_port, S(28) => 
                           routing_wires_7_28_port, S(27) => 
                           routing_wires_7_27_port, S(26) => 
                           routing_wires_7_26_port, S(25) => 
                           routing_wires_7_25_port, S(24) => 
                           routing_wires_7_24_port, S(23) => 
                           routing_wires_7_23_port, S(22) => 
                           routing_wires_7_22_port, S(21) => 
                           routing_wires_7_21_port, S(20) => 
                           routing_wires_7_20_port, S(19) => 
                           routing_wires_7_19_port, S(18) => 
                           routing_wires_7_18_port, S(17) => 
                           routing_wires_7_17_port, S(16) => 
                           routing_wires_7_16_port, S(15) => 
                           routing_wires_7_15_port, S(14) => 
                           routing_wires_7_14_port, S(13) => 
                           routing_wires_7_13_port, S(12) => 
                           routing_wires_7_12_port, S(11) => 
                           routing_wires_7_11_port, S(10) => 
                           routing_wires_7_10_port, S(9) => 
                           routing_wires_7_9_port, S(8) => 
                           routing_wires_7_8_port, S(7) => 
                           routing_wires_7_7_port, S(6) => 
                           routing_wires_7_6_port, S(5) => 
                           routing_wires_7_5_port, S(4) => 
                           routing_wires_7_4_port, S(3) => 
                           routing_wires_7_3_port, S(2) => 
                           routing_wires_7_2_port, S(1) => 
                           routing_wires_7_1_port, S(0) => 
                           routing_wires_7_0_port, Cout => net3148);
   N_shift_pin_port4 <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, 
      n21, n21, n21, n22, n21, n21, n21 );
   gi_8 : generator_N_bit16_4 port map( multiplicant(15) => multiplicand(15), 
      multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin_port4, select_signal(2) => multiplier(9), 
      select_signal(1) => multiplier(8), select_signal(0) => multiplier(7), 
      Out_value(31) => routing_wires_8_31_port, Out_value(30) => 
      routing_wires_8_30_port, Out_value(29) => routing_wires_8_29_port, 
      Out_value(28) => routing_wires_8_28_port, Out_value(27) => 
      routing_wires_8_27_port, Out_value(26) => routing_wires_8_26_port, 
      Out_value(25) => routing_wires_8_25_port, Out_value(24) => 
      routing_wires_8_24_port, Out_value(23) => routing_wires_8_23_port, 
      Out_value(22) => routing_wires_8_22_port, Out_value(21) => 
      routing_wires_8_21_port, Out_value(20) => routing_wires_8_20_port, 
      Out_value(19) => routing_wires_8_19_port, Out_value(18) => 
      routing_wires_8_18_port, Out_value(17) => routing_wires_8_17_port, 
      Out_value(16) => routing_wires_8_16_port, Out_value(15) => 
      routing_wires_8_15_port, Out_value(14) => routing_wires_8_14_port, 
      Out_value(13) => routing_wires_8_13_port, Out_value(12) => 
      routing_wires_8_12_port, Out_value(11) => routing_wires_8_11_port, 
      Out_value(10) => routing_wires_8_10_port, Out_value(9) => 
      routing_wires_8_9_port, Out_value(8) => routing_wires_8_8_port, 
      Out_value(7) => routing_wires_8_7_port, Out_value(6) => 
      routing_wires_8_6_port, Out_value(5) => routing_wires_8_5_port, 
      Out_value(4) => routing_wires_8_4_port, Out_value(3) => 
      routing_wires_8_3_port, Out_value(2) => routing_wires_8_2_port, 
      Out_value(1) => routing_wires_8_1_port, Out_value(0) => 
      routing_wires_8_0_port);
   ai_8 : pentium4_adder_XBIT32_NBIT4_4 port map( A(31) => 
                           routing_wires_7_31_port, A(30) => 
                           routing_wires_7_30_port, A(29) => 
                           routing_wires_7_29_port, A(28) => 
                           routing_wires_7_28_port, A(27) => 
                           routing_wires_7_27_port, A(26) => 
                           routing_wires_7_26_port, A(25) => 
                           routing_wires_7_25_port, A(24) => 
                           routing_wires_7_24_port, A(23) => 
                           routing_wires_7_23_port, A(22) => 
                           routing_wires_7_22_port, A(21) => 
                           routing_wires_7_21_port, A(20) => 
                           routing_wires_7_20_port, A(19) => 
                           routing_wires_7_19_port, A(18) => 
                           routing_wires_7_18_port, A(17) => 
                           routing_wires_7_17_port, A(16) => 
                           routing_wires_7_16_port, A(15) => 
                           routing_wires_7_15_port, A(14) => 
                           routing_wires_7_14_port, A(13) => 
                           routing_wires_7_13_port, A(12) => 
                           routing_wires_7_12_port, A(11) => 
                           routing_wires_7_11_port, A(10) => 
                           routing_wires_7_10_port, A(9) => 
                           routing_wires_7_9_port, A(8) => 
                           routing_wires_7_8_port, A(7) => 
                           routing_wires_7_7_port, A(6) => 
                           routing_wires_7_6_port, A(5) => 
                           routing_wires_7_5_port, A(4) => 
                           routing_wires_7_4_port, A(3) => 
                           routing_wires_7_3_port, A(2) => 
                           routing_wires_7_2_port, A(1) => 
                           routing_wires_7_1_port, A(0) => 
                           routing_wires_7_0_port, B(31) => 
                           routing_wires_8_31_port, B(30) => 
                           routing_wires_8_30_port, B(29) => 
                           routing_wires_8_29_port, B(28) => 
                           routing_wires_8_28_port, B(27) => 
                           routing_wires_8_27_port, B(26) => 
                           routing_wires_8_26_port, B(25) => 
                           routing_wires_8_25_port, B(24) => 
                           routing_wires_8_24_port, B(23) => 
                           routing_wires_8_23_port, B(22) => 
                           routing_wires_8_22_port, B(21) => 
                           routing_wires_8_21_port, B(20) => 
                           routing_wires_8_20_port, B(19) => 
                           routing_wires_8_19_port, B(18) => 
                           routing_wires_8_18_port, B(17) => 
                           routing_wires_8_17_port, B(16) => 
                           routing_wires_8_16_port, B(15) => 
                           routing_wires_8_15_port, B(14) => 
                           routing_wires_8_14_port, B(13) => 
                           routing_wires_8_13_port, B(12) => 
                           routing_wires_8_12_port, B(11) => 
                           routing_wires_8_11_port, B(10) => 
                           routing_wires_8_10_port, B(9) => 
                           routing_wires_8_9_port, B(8) => 
                           routing_wires_8_8_port, B(7) => 
                           routing_wires_8_7_port, B(6) => 
                           routing_wires_8_6_port, B(5) => 
                           routing_wires_8_5_port, B(4) => 
                           routing_wires_8_4_port, B(3) => 
                           routing_wires_8_3_port, B(2) => 
                           routing_wires_8_2_port, B(1) => 
                           routing_wires_8_1_port, B(0) => 
                           routing_wires_8_0_port, C_0 => n21, S(31) => 
                           routing_wires_9_31_port, S(30) => 
                           routing_wires_9_30_port, S(29) => 
                           routing_wires_9_29_port, S(28) => 
                           routing_wires_9_28_port, S(27) => 
                           routing_wires_9_27_port, S(26) => 
                           routing_wires_9_26_port, S(25) => 
                           routing_wires_9_25_port, S(24) => 
                           routing_wires_9_24_port, S(23) => 
                           routing_wires_9_23_port, S(22) => 
                           routing_wires_9_22_port, S(21) => 
                           routing_wires_9_21_port, S(20) => 
                           routing_wires_9_20_port, S(19) => 
                           routing_wires_9_19_port, S(18) => 
                           routing_wires_9_18_port, S(17) => 
                           routing_wires_9_17_port, S(16) => 
                           routing_wires_9_16_port, S(15) => 
                           routing_wires_9_15_port, S(14) => 
                           routing_wires_9_14_port, S(13) => 
                           routing_wires_9_13_port, S(12) => 
                           routing_wires_9_12_port, S(11) => 
                           routing_wires_9_11_port, S(10) => 
                           routing_wires_9_10_port, S(9) => 
                           routing_wires_9_9_port, S(8) => 
                           routing_wires_9_8_port, S(7) => 
                           routing_wires_9_7_port, S(6) => 
                           routing_wires_9_6_port, S(5) => 
                           routing_wires_9_5_port, S(4) => 
                           routing_wires_9_4_port, S(3) => 
                           routing_wires_9_3_port, S(2) => 
                           routing_wires_9_2_port, S(1) => 
                           routing_wires_9_1_port, S(0) => 
                           routing_wires_9_0_port, Cout => net3147);
   N_shift_pin_port5 <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, 
      n21, n21, n21, n22, n21, n22, n21 );
   gi_10 : generator_N_bit16_3 port map( multiplicant(15) => multiplicand(15), 
      multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin_port5, select_signal(2) => multiplier(11), 
      select_signal(1) => multiplier(10), select_signal(0) => multiplier(9), 
      Out_value(31) => routing_wires_10_31_port, Out_value(30) => 
      routing_wires_10_30_port, Out_value(29) => routing_wires_10_29_port, 
      Out_value(28) => routing_wires_10_28_port, Out_value(27) => 
      routing_wires_10_27_port, Out_value(26) => routing_wires_10_26_port, 
      Out_value(25) => routing_wires_10_25_port, Out_value(24) => 
      routing_wires_10_24_port, Out_value(23) => routing_wires_10_23_port, 
      Out_value(22) => routing_wires_10_22_port, Out_value(21) => 
      routing_wires_10_21_port, Out_value(20) => routing_wires_10_20_port, 
      Out_value(19) => routing_wires_10_19_port, Out_value(18) => 
      routing_wires_10_18_port, Out_value(17) => routing_wires_10_17_port, 
      Out_value(16) => routing_wires_10_16_port, Out_value(15) => 
      routing_wires_10_15_port, Out_value(14) => routing_wires_10_14_port, 
      Out_value(13) => routing_wires_10_13_port, Out_value(12) => 
      routing_wires_10_12_port, Out_value(11) => routing_wires_10_11_port, 
      Out_value(10) => routing_wires_10_10_port, Out_value(9) => 
      routing_wires_10_9_port, Out_value(8) => routing_wires_10_8_port, 
      Out_value(7) => routing_wires_10_7_port, Out_value(6) => 
      routing_wires_10_6_port, Out_value(5) => routing_wires_10_5_port, 
      Out_value(4) => routing_wires_10_4_port, Out_value(3) => 
      routing_wires_10_3_port, Out_value(2) => routing_wires_10_2_port, 
      Out_value(1) => routing_wires_10_1_port, Out_value(0) => 
      routing_wires_10_0_port);
   ai_10 : pentium4_adder_XBIT32_NBIT4_3 port map( A(31) => 
                           routing_wires_9_31_port, A(30) => 
                           routing_wires_9_30_port, A(29) => 
                           routing_wires_9_29_port, A(28) => 
                           routing_wires_9_28_port, A(27) => 
                           routing_wires_9_27_port, A(26) => 
                           routing_wires_9_26_port, A(25) => 
                           routing_wires_9_25_port, A(24) => 
                           routing_wires_9_24_port, A(23) => 
                           routing_wires_9_23_port, A(22) => 
                           routing_wires_9_22_port, A(21) => 
                           routing_wires_9_21_port, A(20) => 
                           routing_wires_9_20_port, A(19) => 
                           routing_wires_9_19_port, A(18) => 
                           routing_wires_9_18_port, A(17) => 
                           routing_wires_9_17_port, A(16) => 
                           routing_wires_9_16_port, A(15) => 
                           routing_wires_9_15_port, A(14) => 
                           routing_wires_9_14_port, A(13) => 
                           routing_wires_9_13_port, A(12) => 
                           routing_wires_9_12_port, A(11) => 
                           routing_wires_9_11_port, A(10) => 
                           routing_wires_9_10_port, A(9) => 
                           routing_wires_9_9_port, A(8) => 
                           routing_wires_9_8_port, A(7) => 
                           routing_wires_9_7_port, A(6) => 
                           routing_wires_9_6_port, A(5) => 
                           routing_wires_9_5_port, A(4) => 
                           routing_wires_9_4_port, A(3) => 
                           routing_wires_9_3_port, A(2) => 
                           routing_wires_9_2_port, A(1) => 
                           routing_wires_9_1_port, A(0) => 
                           routing_wires_9_0_port, B(31) => 
                           routing_wires_10_31_port, B(30) => 
                           routing_wires_10_30_port, B(29) => 
                           routing_wires_10_29_port, B(28) => 
                           routing_wires_10_28_port, B(27) => 
                           routing_wires_10_27_port, B(26) => 
                           routing_wires_10_26_port, B(25) => 
                           routing_wires_10_25_port, B(24) => 
                           routing_wires_10_24_port, B(23) => 
                           routing_wires_10_23_port, B(22) => 
                           routing_wires_10_22_port, B(21) => 
                           routing_wires_10_21_port, B(20) => 
                           routing_wires_10_20_port, B(19) => 
                           routing_wires_10_19_port, B(18) => 
                           routing_wires_10_18_port, B(17) => 
                           routing_wires_10_17_port, B(16) => 
                           routing_wires_10_16_port, B(15) => 
                           routing_wires_10_15_port, B(14) => 
                           routing_wires_10_14_port, B(13) => 
                           routing_wires_10_13_port, B(12) => 
                           routing_wires_10_12_port, B(11) => 
                           routing_wires_10_11_port, B(10) => 
                           routing_wires_10_10_port, B(9) => 
                           routing_wires_10_9_port, B(8) => 
                           routing_wires_10_8_port, B(7) => 
                           routing_wires_10_7_port, B(6) => 
                           routing_wires_10_6_port, B(5) => 
                           routing_wires_10_5_port, B(4) => 
                           routing_wires_10_4_port, B(3) => 
                           routing_wires_10_3_port, B(2) => 
                           routing_wires_10_2_port, B(1) => 
                           routing_wires_10_1_port, B(0) => 
                           routing_wires_10_0_port, C_0 => n21, S(31) => 
                           routing_wires_11_31_port, S(30) => 
                           routing_wires_11_30_port, S(29) => 
                           routing_wires_11_29_port, S(28) => 
                           routing_wires_11_28_port, S(27) => 
                           routing_wires_11_27_port, S(26) => 
                           routing_wires_11_26_port, S(25) => 
                           routing_wires_11_25_port, S(24) => 
                           routing_wires_11_24_port, S(23) => 
                           routing_wires_11_23_port, S(22) => 
                           routing_wires_11_22_port, S(21) => 
                           routing_wires_11_21_port, S(20) => 
                           routing_wires_11_20_port, S(19) => 
                           routing_wires_11_19_port, S(18) => 
                           routing_wires_11_18_port, S(17) => 
                           routing_wires_11_17_port, S(16) => 
                           routing_wires_11_16_port, S(15) => 
                           routing_wires_11_15_port, S(14) => 
                           routing_wires_11_14_port, S(13) => 
                           routing_wires_11_13_port, S(12) => 
                           routing_wires_11_12_port, S(11) => 
                           routing_wires_11_11_port, S(10) => 
                           routing_wires_11_10_port, S(9) => 
                           routing_wires_11_9_port, S(8) => 
                           routing_wires_11_8_port, S(7) => 
                           routing_wires_11_7_port, S(6) => 
                           routing_wires_11_6_port, S(5) => 
                           routing_wires_11_5_port, S(4) => 
                           routing_wires_11_4_port, S(3) => 
                           routing_wires_11_3_port, S(2) => 
                           routing_wires_11_2_port, S(1) => 
                           routing_wires_11_1_port, S(0) => 
                           routing_wires_11_0_port, Cout => net3146);
   N_shift_pin_port6 <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, 
      n21, n21, n21, n22, n22, n21, n21 );
   gi_12 : generator_N_bit16_2 port map( multiplicant(15) => multiplicand(15), 
      multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin_port6, select_signal(2) => multiplier(13), 
      select_signal(1) => multiplier(12), select_signal(0) => multiplier(11), 
      Out_value(31) => routing_wires_12_31_port, Out_value(30) => 
      routing_wires_12_30_port, Out_value(29) => routing_wires_12_29_port, 
      Out_value(28) => routing_wires_12_28_port, Out_value(27) => 
      routing_wires_12_27_port, Out_value(26) => routing_wires_12_26_port, 
      Out_value(25) => routing_wires_12_25_port, Out_value(24) => 
      routing_wires_12_24_port, Out_value(23) => routing_wires_12_23_port, 
      Out_value(22) => routing_wires_12_22_port, Out_value(21) => 
      routing_wires_12_21_port, Out_value(20) => routing_wires_12_20_port, 
      Out_value(19) => routing_wires_12_19_port, Out_value(18) => 
      routing_wires_12_18_port, Out_value(17) => routing_wires_12_17_port, 
      Out_value(16) => routing_wires_12_16_port, Out_value(15) => 
      routing_wires_12_15_port, Out_value(14) => routing_wires_12_14_port, 
      Out_value(13) => routing_wires_12_13_port, Out_value(12) => 
      routing_wires_12_12_port, Out_value(11) => routing_wires_12_11_port, 
      Out_value(10) => routing_wires_12_10_port, Out_value(9) => 
      routing_wires_12_9_port, Out_value(8) => routing_wires_12_8_port, 
      Out_value(7) => routing_wires_12_7_port, Out_value(6) => 
      routing_wires_12_6_port, Out_value(5) => routing_wires_12_5_port, 
      Out_value(4) => routing_wires_12_4_port, Out_value(3) => 
      routing_wires_12_3_port, Out_value(2) => routing_wires_12_2_port, 
      Out_value(1) => routing_wires_12_1_port, Out_value(0) => 
      routing_wires_12_0_port);
   ai_12 : pentium4_adder_XBIT32_NBIT4_2 port map( A(31) => 
                           routing_wires_11_31_port, A(30) => 
                           routing_wires_11_30_port, A(29) => 
                           routing_wires_11_29_port, A(28) => 
                           routing_wires_11_28_port, A(27) => 
                           routing_wires_11_27_port, A(26) => 
                           routing_wires_11_26_port, A(25) => 
                           routing_wires_11_25_port, A(24) => 
                           routing_wires_11_24_port, A(23) => 
                           routing_wires_11_23_port, A(22) => 
                           routing_wires_11_22_port, A(21) => 
                           routing_wires_11_21_port, A(20) => 
                           routing_wires_11_20_port, A(19) => 
                           routing_wires_11_19_port, A(18) => 
                           routing_wires_11_18_port, A(17) => 
                           routing_wires_11_17_port, A(16) => 
                           routing_wires_11_16_port, A(15) => 
                           routing_wires_11_15_port, A(14) => 
                           routing_wires_11_14_port, A(13) => 
                           routing_wires_11_13_port, A(12) => 
                           routing_wires_11_12_port, A(11) => 
                           routing_wires_11_11_port, A(10) => 
                           routing_wires_11_10_port, A(9) => 
                           routing_wires_11_9_port, A(8) => 
                           routing_wires_11_8_port, A(7) => 
                           routing_wires_11_7_port, A(6) => 
                           routing_wires_11_6_port, A(5) => 
                           routing_wires_11_5_port, A(4) => 
                           routing_wires_11_4_port, A(3) => 
                           routing_wires_11_3_port, A(2) => 
                           routing_wires_11_2_port, A(1) => 
                           routing_wires_11_1_port, A(0) => 
                           routing_wires_11_0_port, B(31) => 
                           routing_wires_12_31_port, B(30) => 
                           routing_wires_12_30_port, B(29) => 
                           routing_wires_12_29_port, B(28) => 
                           routing_wires_12_28_port, B(27) => 
                           routing_wires_12_27_port, B(26) => 
                           routing_wires_12_26_port, B(25) => 
                           routing_wires_12_25_port, B(24) => 
                           routing_wires_12_24_port, B(23) => 
                           routing_wires_12_23_port, B(22) => 
                           routing_wires_12_22_port, B(21) => 
                           routing_wires_12_21_port, B(20) => 
                           routing_wires_12_20_port, B(19) => 
                           routing_wires_12_19_port, B(18) => 
                           routing_wires_12_18_port, B(17) => 
                           routing_wires_12_17_port, B(16) => 
                           routing_wires_12_16_port, B(15) => 
                           routing_wires_12_15_port, B(14) => 
                           routing_wires_12_14_port, B(13) => 
                           routing_wires_12_13_port, B(12) => 
                           routing_wires_12_12_port, B(11) => 
                           routing_wires_12_11_port, B(10) => 
                           routing_wires_12_10_port, B(9) => 
                           routing_wires_12_9_port, B(8) => 
                           routing_wires_12_8_port, B(7) => 
                           routing_wires_12_7_port, B(6) => 
                           routing_wires_12_6_port, B(5) => 
                           routing_wires_12_5_port, B(4) => 
                           routing_wires_12_4_port, B(3) => 
                           routing_wires_12_3_port, B(2) => 
                           routing_wires_12_2_port, B(1) => 
                           routing_wires_12_1_port, B(0) => 
                           routing_wires_12_0_port, C_0 => n21, S(31) => 
                           routing_wires_13_31_port, S(30) => 
                           routing_wires_13_30_port, S(29) => 
                           routing_wires_13_29_port, S(28) => 
                           routing_wires_13_28_port, S(27) => 
                           routing_wires_13_27_port, S(26) => 
                           routing_wires_13_26_port, S(25) => 
                           routing_wires_13_25_port, S(24) => 
                           routing_wires_13_24_port, S(23) => 
                           routing_wires_13_23_port, S(22) => 
                           routing_wires_13_22_port, S(21) => 
                           routing_wires_13_21_port, S(20) => 
                           routing_wires_13_20_port, S(19) => 
                           routing_wires_13_19_port, S(18) => 
                           routing_wires_13_18_port, S(17) => 
                           routing_wires_13_17_port, S(16) => 
                           routing_wires_13_16_port, S(15) => 
                           routing_wires_13_15_port, S(14) => 
                           routing_wires_13_14_port, S(13) => 
                           routing_wires_13_13_port, S(12) => 
                           routing_wires_13_12_port, S(11) => 
                           routing_wires_13_11_port, S(10) => 
                           routing_wires_13_10_port, S(9) => 
                           routing_wires_13_9_port, S(8) => 
                           routing_wires_13_8_port, S(7) => 
                           routing_wires_13_7_port, S(6) => 
                           routing_wires_13_6_port, S(5) => 
                           routing_wires_13_5_port, S(4) => 
                           routing_wires_13_4_port, S(3) => 
                           routing_wires_13_3_port, S(2) => 
                           routing_wires_13_2_port, S(1) => 
                           routing_wires_13_1_port, S(0) => 
                           routing_wires_13_0_port, Cout => net3145);
   N_shift_pin_port7 <= ( n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21
      , n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, n21, 
      n21, n21, n21, n22, n22, n22, n21 );
   gi_l_14 : generator_N_bit16_1 port map( multiplicant(15) => multiplicand(15)
      , multiplicant(14) => multiplicand(14), multiplicant(13) => 
      multiplicand(13), multiplicant(12) => multiplicand(12), multiplicant(11) 
      => multiplicand(11), multiplicant(10) => multiplicand(10), 
      multiplicant(9) => multiplicand(9), multiplicant(8) => multiplicand(8), 
      multiplicant(7) => multiplicand(7), multiplicant(6) => multiplicand(6), 
      multiplicant(5) => multiplicand(5), multiplicant(4) => multiplicand(4), 
      multiplicant(3) => multiplicand(3), multiplicant(2) => multiplicand(2), 
      multiplicant(1) => multiplicand(1), multiplicant(0) => multiplicand(0), 
      N_shift => N_shift_pin_port7, select_signal(2) => multiplier(15), 
      select_signal(1) => multiplier(14), select_signal(0) => multiplier(13), 
      Out_value(31) => routing_wires_14_31_port, Out_value(30) => 
      routing_wires_14_30_port, Out_value(29) => routing_wires_14_29_port, 
      Out_value(28) => routing_wires_14_28_port, Out_value(27) => 
      routing_wires_14_27_port, Out_value(26) => routing_wires_14_26_port, 
      Out_value(25) => routing_wires_14_25_port, Out_value(24) => 
      routing_wires_14_24_port, Out_value(23) => routing_wires_14_23_port, 
      Out_value(22) => routing_wires_14_22_port, Out_value(21) => 
      routing_wires_14_21_port, Out_value(20) => routing_wires_14_20_port, 
      Out_value(19) => routing_wires_14_19_port, Out_value(18) => 
      routing_wires_14_18_port, Out_value(17) => routing_wires_14_17_port, 
      Out_value(16) => routing_wires_14_16_port, Out_value(15) => 
      routing_wires_14_15_port, Out_value(14) => routing_wires_14_14_port, 
      Out_value(13) => routing_wires_14_13_port, Out_value(12) => 
      routing_wires_14_12_port, Out_value(11) => routing_wires_14_11_port, 
      Out_value(10) => routing_wires_14_10_port, Out_value(9) => 
      routing_wires_14_9_port, Out_value(8) => routing_wires_14_8_port, 
      Out_value(7) => routing_wires_14_7_port, Out_value(6) => 
      routing_wires_14_6_port, Out_value(5) => routing_wires_14_5_port, 
      Out_value(4) => routing_wires_14_4_port, Out_value(3) => 
      routing_wires_14_3_port, Out_value(2) => routing_wires_14_2_port, 
      Out_value(1) => routing_wires_14_1_port, Out_value(0) => 
      routing_wires_14_0_port);
   ai_l_14 : pentium4_adder_XBIT32_NBIT4_1 port map( A(31) => 
                           routing_wires_13_31_port, A(30) => 
                           routing_wires_13_30_port, A(29) => 
                           routing_wires_13_29_port, A(28) => 
                           routing_wires_13_28_port, A(27) => 
                           routing_wires_13_27_port, A(26) => 
                           routing_wires_13_26_port, A(25) => 
                           routing_wires_13_25_port, A(24) => 
                           routing_wires_13_24_port, A(23) => 
                           routing_wires_13_23_port, A(22) => 
                           routing_wires_13_22_port, A(21) => 
                           routing_wires_13_21_port, A(20) => 
                           routing_wires_13_20_port, A(19) => 
                           routing_wires_13_19_port, A(18) => 
                           routing_wires_13_18_port, A(17) => 
                           routing_wires_13_17_port, A(16) => 
                           routing_wires_13_16_port, A(15) => 
                           routing_wires_13_15_port, A(14) => 
                           routing_wires_13_14_port, A(13) => 
                           routing_wires_13_13_port, A(12) => 
                           routing_wires_13_12_port, A(11) => 
                           routing_wires_13_11_port, A(10) => 
                           routing_wires_13_10_port, A(9) => 
                           routing_wires_13_9_port, A(8) => 
                           routing_wires_13_8_port, A(7) => 
                           routing_wires_13_7_port, A(6) => 
                           routing_wires_13_6_port, A(5) => 
                           routing_wires_13_5_port, A(4) => 
                           routing_wires_13_4_port, A(3) => 
                           routing_wires_13_3_port, A(2) => 
                           routing_wires_13_2_port, A(1) => 
                           routing_wires_13_1_port, A(0) => 
                           routing_wires_13_0_port, B(31) => 
                           routing_wires_14_31_port, B(30) => 
                           routing_wires_14_30_port, B(29) => 
                           routing_wires_14_29_port, B(28) => 
                           routing_wires_14_28_port, B(27) => 
                           routing_wires_14_27_port, B(26) => 
                           routing_wires_14_26_port, B(25) => 
                           routing_wires_14_25_port, B(24) => 
                           routing_wires_14_24_port, B(23) => 
                           routing_wires_14_23_port, B(22) => 
                           routing_wires_14_22_port, B(21) => 
                           routing_wires_14_21_port, B(20) => 
                           routing_wires_14_20_port, B(19) => 
                           routing_wires_14_19_port, B(18) => 
                           routing_wires_14_18_port, B(17) => 
                           routing_wires_14_17_port, B(16) => 
                           routing_wires_14_16_port, B(15) => 
                           routing_wires_14_15_port, B(14) => 
                           routing_wires_14_14_port, B(13) => 
                           routing_wires_14_13_port, B(12) => 
                           routing_wires_14_12_port, B(11) => 
                           routing_wires_14_11_port, B(10) => 
                           routing_wires_14_10_port, B(9) => 
                           routing_wires_14_9_port, B(8) => 
                           routing_wires_14_8_port, B(7) => 
                           routing_wires_14_7_port, B(6) => 
                           routing_wires_14_6_port, B(5) => 
                           routing_wires_14_5_port, B(4) => 
                           routing_wires_14_4_port, B(3) => 
                           routing_wires_14_3_port, B(2) => 
                           routing_wires_14_2_port, B(1) => 
                           routing_wires_14_1_port, B(0) => 
                           routing_wires_14_0_port, C_0 => n21, S(31) => 
                           product(31), S(30) => product(30), S(29) => 
                           product(29), S(28) => product(28), S(27) => 
                           product(27), S(26) => product(26), S(25) => 
                           product(25), S(24) => product(24), S(23) => 
                           product(23), S(22) => product(22), S(21) => 
                           product(21), S(20) => product(20), S(19) => 
                           product(19), S(18) => product(18), S(17) => 
                           product(17), S(16) => product(16), S(15) => 
                           product(15), S(14) => product(14), S(13) => 
                           product(13), S(12) => product(12), S(11) => 
                           product(11), S(10) => product(10), S(9) => 
                           product(9), S(8) => product(8), S(7) => product(7), 
                           S(6) => product(6), S(5) => product(5), S(4) => 
                           product(4), S(3) => product(3), S(2) => product(2), 
                           S(1) => product(1), S(0) => product(0), Cout => 
                           net3144);
   n21 <= '0';
   n22 <= '1';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity Shifter_NBIT32 is

   port( left_right, logic_Arith, shift_rot : in std_logic;  a, b : in 
         std_logic_vector (31 downto 0);  o : out std_logic_vector (31 downto 
         0));

end Shifter_NBIT32;

architecture SYN_beh of Shifter_NBIT32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Shifter_NBIT32_DW_rbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_NBIT32_DW_lbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_NBIT32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_NBIT32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component Shifter_NBIT32_DW_sla_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_NBIT32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   signal N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, 
      N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37
      , N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, 
      N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66
      , N67, N68, N69, N70, N71, N72, N108, N109, N110, N111, N112, N113, N114,
      N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, 
      N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, 
      N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, 
      N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, 
      N163, N164, N165, N166, N167, N168, N169, N170, N171, N205, N206, N207, 
      N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, 
      N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, 
      N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, 
      N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, 
      N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
      N268, n7, n8, n9_port, n10_port, n11_port, n12_port, n16_port, n17_port, 
      n18_port, n19_port, n20_port, n21_port, n22_port, n23_port, n24_port, 
      n25_port, n26_port, n27_port, n28_port, n29_port, n30_port, n31_port, 
      n32_port, n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, 
      n39_port, n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, 
      n46_port, n47_port, n48_port, n49_port, n50_port, n51_port, n52_port, 
      n53_port, n54_port, n55_port, n56_port, n57_port, n58_port, n59_port, 
      n60_port, n61_port, n62_port, n63_port, n64_port, n65_port, n66_port, 
      n67_port, n68_port, n69_port, n70_port, n71_port, n72_port, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n206_port, n207_port, n208_port, n209_port, n210_port, n211_port, 
      n212_port, n213_port, n214_port, n215_port, n216_port, n217_port, 
      n218_port, n219_port, n220_port, n221_port, n222_port, n223_port, 
      n224_port, n225_port : std_logic;

begin
   
   n7 <= '0';
   n8 <= '0';
   n9_port <= '0';
   n10_port <= '0';
   n11_port <= '0';
   n12_port <= '0';
   C93 : Shifter_NBIT32_DW01_ash_0 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), DATA_TC => n10_port, SH(4) => 
                           n225_port, SH(3) => n224_port, SH(2) => b(2), SH(1) 
                           => b(1), SH(0) => b(0), SH_TC => n10_port, B(31) => 
                           N268, B(30) => N267, B(29) => N266, B(28) => N265, 
                           B(27) => N264, B(26) => N263, B(25) => N262, B(24) 
                           => N261, B(23) => N260, B(22) => N259, B(21) => N258
                           , B(20) => N257, B(19) => N256, B(18) => N255, B(17)
                           => N254, B(16) => N253, B(15) => N252, B(14) => N251
                           , B(13) => N250, B(12) => N249, B(11) => N248, B(10)
                           => N247, B(9) => N246, B(8) => N245, B(7) => N244, 
                           B(6) => N243, B(5) => N242, B(4) => N241, B(3) => 
                           N240, B(2) => N239, B(1) => N238, B(0) => N237);
   C91 : Shifter_NBIT32_DW_sla_0 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n225_port, SH(3) => 
                           n224_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n11_port, B(31) => N236, B(30) => 
                           N235, B(29) => N234, B(28) => N233, B(27) => N232, 
                           B(26) => N231, B(25) => N230, B(24) => N229, B(23) 
                           => N228, B(22) => N227, B(21) => N226, B(20) => N225
                           , B(19) => N224, B(18) => N223, B(17) => N222, B(16)
                           => N221, B(15) => N220, B(14) => N219, B(13) => N218
                           , B(12) => N217, B(11) => N216, B(10) => N215, B(9) 
                           => N214, B(8) => N213, B(7) => N212, B(6) => N211, 
                           B(5) => N210, B(4) => N209, B(3) => N208, B(2) => 
                           N207, B(1) => N206, B(0) => N205);
   C54 : Shifter_NBIT32_DW_rash_0 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), DATA_TC => n12_port, SH(4) => 
                           n225_port, SH(3) => n224_port, SH(2) => b(2), SH(1) 
                           => b(1), SH(0) => b(0), SH_TC => n12_port, B(31) => 
                           N171, B(30) => N170, B(29) => N169, B(28) => N168, 
                           B(27) => N167, B(26) => N166, B(25) => N165, B(24) 
                           => N164, B(23) => N163, B(22) => N162, B(21) => N161
                           , B(20) => N160, B(19) => N159, B(18) => N158, B(17)
                           => N157, B(16) => N156, B(15) => N155, B(14) => N154
                           , B(13) => N153, B(12) => N152, B(11) => N151, B(10)
                           => N150, B(9) => N149, B(8) => N148, B(7) => N147, 
                           B(6) => N146, B(5) => N145, B(4) => N144, B(3) => 
                           N143, B(2) => N142, B(1) => N141, B(0) => N140);
   C52 : Shifter_NBIT32_DW_sra_0 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n225_port, SH(3) => 
                           n224_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n7, B(31) => N139, B(30) => N138, 
                           B(29) => N137, B(28) => N136, B(27) => N135, B(26) 
                           => N134, B(25) => N133, B(24) => N132, B(23) => N131
                           , B(22) => N130, B(21) => N129, B(20) => N128, B(19)
                           => N127, B(18) => N126, B(17) => N125, B(16) => N124
                           , B(15) => N123, B(14) => N122, B(13) => N121, B(12)
                           => N120, B(11) => N119, B(10) => N118, B(9) => N117,
                           B(8) => N116, B(7) => N115, B(6) => N114, B(5) => 
                           N113, B(4) => N112, B(3) => N111, B(2) => N110, B(1)
                           => N109, B(0) => N108);
   C12 : Shifter_NBIT32_DW_lbsh_0 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n225_port, SH(3) => 
                           n224_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n8, B(31) => N72, B(30) => N71, B(29)
                           => N70, B(28) => N69, B(27) => N68, B(26) => N67, 
                           B(25) => N66, B(24) => N65, B(23) => N64, B(22) => 
                           N63, B(21) => N62, B(20) => N61, B(19) => N60, B(18)
                           => N59, B(17) => N58, B(16) => N57, B(15) => N56, 
                           B(14) => N55, B(13) => N54, B(12) => N53, B(11) => 
                           N52, B(10) => N51, B(9) => N50, B(8) => N49, B(7) =>
                           N48, B(6) => N47, B(5) => N46, B(4) => N45, B(3) => 
                           N44, B(2) => N43, B(1) => N42, B(0) => N41);
   C10 : Shifter_NBIT32_DW_rbsh_0 port map( A(31) => a(31), A(30) => a(30), 
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n225_port, SH(3) => 
                           n224_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n9_port, B(31) => N40, B(30) => N39, 
                           B(29) => N38, B(28) => N37, B(27) => N36, B(26) => 
                           N35, B(25) => N34, B(24) => N33, B(23) => N32, B(22)
                           => N31, B(21) => N30, B(20) => N29, B(19) => N28, 
                           B(18) => N27, B(17) => N26, B(16) => N25, B(15) => 
                           N24, B(14) => N23, B(13) => N22, B(12) => N21, B(11)
                           => N20, B(10) => N19, B(9) => N18, B(8) => N17, B(7)
                           => N16, B(6) => N15, B(5) => N14, B(4) => N13, B(3) 
                           => N12, B(2) => N11, B(1) => N10, B(0) => N9);
   U5 : BUF_X1 port map( A => b(3), Z => n224_port);
   U6 : BUF_X1 port map( A => n21_port, Z => n213_port);
   U7 : BUF_X1 port map( A => n21_port, Z => n212_port);
   U8 : BUF_X1 port map( A => n21_port, Z => n214_port);
   U9 : BUF_X1 port map( A => n22_port, Z => n210_port);
   U10 : BUF_X1 port map( A => n22_port, Z => n209_port);
   U13 : NOR2_X1 port map( A1 => n88, A2 => n87, ZN => n21_port);
   U14 : BUF_X1 port map( A => n20_port, Z => n216_port);
   U15 : BUF_X1 port map( A => n20_port, Z => n215_port);
   U16 : BUF_X1 port map( A => n23_port, Z => n207_port);
   U17 : BUF_X1 port map( A => n23_port, Z => n206_port);
   U18 : BUF_X1 port map( A => n22_port, Z => n211_port);
   U19 : BUF_X1 port map( A => n20_port, Z => n217_port);
   U20 : BUF_X1 port map( A => n23_port, Z => n208_port);
   U21 : NOR3_X1 port map( A1 => left_right, A2 => shift_rot, A3 => n86, ZN => 
                           n20_port);
   U22 : NOR3_X1 port map( A1 => n86, A2 => shift_rot, A3 => n87, ZN => 
                           n22_port);
   U23 : AOI222_X1 port map( A1 => N18, A2 => n214_port, B1 => N117, B2 => 
                           n211_port, C1 => N50, C2 => n208_port, ZN => 
                           n16_port);
   U24 : AOI222_X1 port map( A1 => N17, A2 => n214_port, B1 => N116, B2 => 
                           n211_port, C1 => N49, C2 => n208_port, ZN => 
                           n24_port);
   U25 : AOI222_X1 port map( A1 => N22, A2 => n212_port, B1 => N121, B2 => 
                           n209_port, C1 => N54, C2 => n206_port, ZN => n76);
   U26 : AOI222_X1 port map( A1 => N21, A2 => n212_port, B1 => N120, B2 => 
                           n209_port, C1 => N53, C2 => n206_port, ZN => n78);
   U27 : AOI222_X1 port map( A1 => N20, A2 => n212_port, B1 => N119, B2 => 
                           n209_port, C1 => N52, C2 => n206_port, ZN => n80);
   U28 : AOI222_X1 port map( A1 => N19, A2 => n212_port, B1 => N118, B2 => 
                           n209_port, C1 => N51, C2 => n206_port, ZN => n82);
   U29 : BUF_X1 port map( A => n18_port, Z => n222_port);
   U30 : BUF_X1 port map( A => n18_port, Z => n221_port);
   U31 : BUF_X1 port map( A => n19_port, Z => n219_port);
   U32 : BUF_X1 port map( A => n19_port, Z => n218_port);
   U33 : NOR2_X1 port map( A1 => n88, A2 => left_right, ZN => n23_port);
   U34 : BUF_X1 port map( A => n19_port, Z => n220_port);
   U35 : BUF_X1 port map( A => n18_port, Z => n223_port);
   U36 : INV_X1 port map( A => shift_rot, ZN => n88);
   U37 : INV_X1 port map( A => left_right, ZN => n87);
   U38 : AOI222_X1 port map( A1 => N149, A2 => n223_port, B1 => N246, B2 => 
                           n220_port, C1 => N214, C2 => n217_port, ZN => 
                           n17_port);
   U39 : AOI222_X1 port map( A1 => N148, A2 => n223_port, B1 => N245, B2 => 
                           n220_port, C1 => N213, C2 => n217_port, ZN => 
                           n25_port);
   U40 : AOI222_X1 port map( A1 => N147, A2 => n223_port, B1 => N244, B2 => 
                           n220_port, C1 => N212, C2 => n217_port, ZN => 
                           n27_port);
   U41 : AOI222_X1 port map( A1 => N146, A2 => n223_port, B1 => N243, B2 => 
                           n220_port, C1 => N211, C2 => n217_port, ZN => 
                           n29_port);
   U42 : AOI222_X1 port map( A1 => N145, A2 => n223_port, B1 => N242, B2 => 
                           n220_port, C1 => N210, C2 => n217_port, ZN => 
                           n31_port);
   U43 : AOI222_X1 port map( A1 => N144, A2 => n223_port, B1 => N241, B2 => 
                           n220_port, C1 => N209, C2 => n217_port, ZN => 
                           n33_port);
   U44 : AOI222_X1 port map( A1 => N143, A2 => n223_port, B1 => N240, B2 => 
                           n220_port, C1 => N208, C2 => n217_port, ZN => 
                           n35_port);
   U45 : AOI222_X1 port map( A1 => N171, A2 => n223_port, B1 => N268, B2 => 
                           n220_port, C1 => N236, C2 => n217_port, ZN => 
                           n37_port);
   U46 : AOI222_X1 port map( A1 => N155, A2 => n221_port, B1 => N252, B2 => 
                           n218_port, C1 => N220, C2 => n215_port, ZN => n73);
   U47 : AOI222_X1 port map( A1 => N154, A2 => n221_port, B1 => N251, B2 => 
                           n218_port, C1 => N219, C2 => n215_port, ZN => n75);
   U48 : AOI222_X1 port map( A1 => N153, A2 => n221_port, B1 => N250, B2 => 
                           n218_port, C1 => N218, C2 => n215_port, ZN => n77);
   U49 : AOI222_X1 port map( A1 => N152, A2 => n221_port, B1 => N249, B2 => 
                           n218_port, C1 => N217, C2 => n215_port, ZN => n79);
   U50 : AOI222_X1 port map( A1 => N151, A2 => n221_port, B1 => N248, B2 => 
                           n218_port, C1 => N216, C2 => n215_port, ZN => n81);
   U51 : AOI222_X1 port map( A1 => N150, A2 => n221_port, B1 => N247, B2 => 
                           n218_port, C1 => N215, C2 => n215_port, ZN => n83);
   U52 : AOI222_X1 port map( A1 => N142, A2 => n222_port, B1 => N239, B2 => 
                           n219_port, C1 => N207, C2 => n216_port, ZN => 
                           n41_port);
   U53 : AOI222_X1 port map( A1 => N141, A2 => n221_port, B1 => N238, B2 => 
                           n218_port, C1 => N206, C2 => n215_port, ZN => 
                           n63_port);
   U54 : AOI222_X1 port map( A1 => N170, A2 => n222_port, B1 => N267, B2 => 
                           n219_port, C1 => N235, C2 => n216_port, ZN => 
                           n39_port);
   U55 : AOI222_X1 port map( A1 => N169, A2 => n222_port, B1 => N266, B2 => 
                           n219_port, C1 => N234, C2 => n216_port, ZN => 
                           n43_port);
   U56 : AOI222_X1 port map( A1 => N168, A2 => n222_port, B1 => N265, B2 => 
                           n219_port, C1 => N233, C2 => n216_port, ZN => 
                           n45_port);
   U57 : AOI222_X1 port map( A1 => N167, A2 => n222_port, B1 => N264, B2 => 
                           n219_port, C1 => N232, C2 => n216_port, ZN => 
                           n47_port);
   U58 : AOI222_X1 port map( A1 => N166, A2 => n222_port, B1 => N263, B2 => 
                           n219_port, C1 => N231, C2 => n216_port, ZN => 
                           n49_port);
   U59 : AOI222_X1 port map( A1 => N165, A2 => n222_port, B1 => N262, B2 => 
                           n219_port, C1 => N230, C2 => n216_port, ZN => 
                           n51_port);
   U60 : AOI222_X1 port map( A1 => N164, A2 => n222_port, B1 => N261, B2 => 
                           n219_port, C1 => N229, C2 => n216_port, ZN => 
                           n53_port);
   U61 : AOI222_X1 port map( A1 => N163, A2 => n222_port, B1 => N260, B2 => 
                           n219_port, C1 => N228, C2 => n216_port, ZN => 
                           n55_port);
   U62 : AOI222_X1 port map( A1 => N162, A2 => n222_port, B1 => N259, B2 => 
                           n219_port, C1 => N227, C2 => n216_port, ZN => 
                           n57_port);
   U63 : AOI222_X1 port map( A1 => N161, A2 => n222_port, B1 => N258, B2 => 
                           n219_port, C1 => N226, C2 => n216_port, ZN => 
                           n59_port);
   U64 : AOI222_X1 port map( A1 => N160, A2 => n222_port, B1 => N257, B2 => 
                           n219_port, C1 => N225, C2 => n216_port, ZN => 
                           n61_port);
   U65 : AOI222_X1 port map( A1 => N159, A2 => n221_port, B1 => N256, B2 => 
                           n218_port, C1 => N224, C2 => n215_port, ZN => 
                           n65_port);
   U66 : AOI222_X1 port map( A1 => N158, A2 => n221_port, B1 => N255, B2 => 
                           n218_port, C1 => N223, C2 => n215_port, ZN => 
                           n67_port);
   U67 : AOI222_X1 port map( A1 => N157, A2 => n221_port, B1 => N254, B2 => 
                           n218_port, C1 => N222, C2 => n215_port, ZN => 
                           n69_port);
   U68 : AOI222_X1 port map( A1 => N156, A2 => n221_port, B1 => N253, B2 => 
                           n218_port, C1 => N221, C2 => n215_port, ZN => 
                           n71_port);
   U69 : NOR3_X1 port map( A1 => logic_Arith, A2 => shift_rot, A3 => left_right
                           , ZN => n19_port);
   U70 : AOI222_X1 port map( A1 => N16, A2 => n214_port, B1 => N115, B2 => 
                           n211_port, C1 => N48, C2 => n208_port, ZN => 
                           n26_port);
   U71 : AOI222_X1 port map( A1 => N15, A2 => n214_port, B1 => N114, B2 => 
                           n211_port, C1 => N47, C2 => n208_port, ZN => 
                           n28_port);
   U72 : AOI222_X1 port map( A1 => N14, A2 => n214_port, B1 => N113, B2 => 
                           n211_port, C1 => N46, C2 => n208_port, ZN => 
                           n30_port);
   U73 : AOI222_X1 port map( A1 => N13, A2 => n214_port, B1 => N112, B2 => 
                           n211_port, C1 => N45, C2 => n208_port, ZN => 
                           n32_port);
   U74 : AOI222_X1 port map( A1 => N12, A2 => n214_port, B1 => N111, B2 => 
                           n211_port, C1 => N44, C2 => n208_port, ZN => 
                           n34_port);
   U75 : AOI222_X1 port map( A1 => N24, A2 => n212_port, B1 => N123, B2 => 
                           n209_port, C1 => N56, C2 => n206_port, ZN => 
                           n72_port);
   U76 : AOI222_X1 port map( A1 => N23, A2 => n212_port, B1 => N122, B2 => 
                           n209_port, C1 => N55, C2 => n206_port, ZN => n74);
   U77 : AOI222_X1 port map( A1 => N11, A2 => n213_port, B1 => N110, B2 => 
                           n210_port, C1 => N43, C2 => n207_port, ZN => 
                           n40_port);
   U78 : AOI222_X1 port map( A1 => N10, A2 => n212_port, B1 => N109, B2 => 
                           n209_port, C1 => N42, C2 => n206_port, ZN => 
                           n62_port);
   U79 : AOI222_X1 port map( A1 => N9, A2 => n212_port, B1 => N108, B2 => 
                           n209_port, C1 => N41, C2 => n206_port, ZN => n84);
   U80 : AOI222_X1 port map( A1 => N39, A2 => n213_port, B1 => N138, B2 => 
                           n210_port, C1 => N71, C2 => n207_port, ZN => 
                           n38_port);
   U81 : AOI222_X1 port map( A1 => N38, A2 => n213_port, B1 => N137, B2 => 
                           n210_port, C1 => N70, C2 => n207_port, ZN => 
                           n42_port);
   U82 : AOI222_X1 port map( A1 => N37, A2 => n213_port, B1 => N136, B2 => 
                           n210_port, C1 => N69, C2 => n207_port, ZN => 
                           n44_port);
   U83 : AOI222_X1 port map( A1 => N36, A2 => n213_port, B1 => N135, B2 => 
                           n210_port, C1 => N68, C2 => n207_port, ZN => 
                           n46_port);
   U84 : AOI222_X1 port map( A1 => N35, A2 => n213_port, B1 => N134, B2 => 
                           n210_port, C1 => N67, C2 => n207_port, ZN => 
                           n48_port);
   U85 : AOI222_X1 port map( A1 => N34, A2 => n213_port, B1 => N133, B2 => 
                           n210_port, C1 => N66, C2 => n207_port, ZN => 
                           n50_port);
   U86 : AOI222_X1 port map( A1 => N33, A2 => n213_port, B1 => N132, B2 => 
                           n210_port, C1 => N65, C2 => n207_port, ZN => 
                           n52_port);
   U87 : AOI222_X1 port map( A1 => N32, A2 => n213_port, B1 => N131, B2 => 
                           n210_port, C1 => N64, C2 => n207_port, ZN => 
                           n54_port);
   U88 : AOI222_X1 port map( A1 => N31, A2 => n213_port, B1 => N130, B2 => 
                           n210_port, C1 => N63, C2 => n207_port, ZN => 
                           n56_port);
   U89 : AOI222_X1 port map( A1 => N30, A2 => n213_port, B1 => N129, B2 => 
                           n210_port, C1 => N62, C2 => n207_port, ZN => 
                           n58_port);
   U90 : AOI222_X1 port map( A1 => N29, A2 => n213_port, B1 => N128, B2 => 
                           n210_port, C1 => N61, C2 => n207_port, ZN => 
                           n60_port);
   U91 : AOI222_X1 port map( A1 => N28, A2 => n212_port, B1 => N127, B2 => 
                           n209_port, C1 => N60, C2 => n206_port, ZN => 
                           n64_port);
   U92 : AOI222_X1 port map( A1 => N27, A2 => n212_port, B1 => N126, B2 => 
                           n209_port, C1 => N59, C2 => n206_port, ZN => 
                           n66_port);
   U93 : AOI222_X1 port map( A1 => N26, A2 => n212_port, B1 => N125, B2 => 
                           n209_port, C1 => N58, C2 => n206_port, ZN => 
                           n68_port);
   U94 : AOI222_X1 port map( A1 => N25, A2 => n212_port, B1 => N124, B2 => 
                           n209_port, C1 => N57, C2 => n206_port, ZN => 
                           n70_port);
   U95 : NOR3_X1 port map( A1 => logic_Arith, A2 => shift_rot, A3 => n87, ZN =>
                           n18_port);
   U96 : INV_X1 port map( A => logic_Arith, ZN => n86);
   U97 : AOI222_X1 port map( A1 => N140, A2 => n221_port, B1 => N237, B2 => 
                           n218_port, C1 => N205, C2 => n215_port, ZN => n85);
   U98 : AOI222_X1 port map( A1 => N40, A2 => n214_port, B1 => N139, B2 => 
                           n211_port, C1 => N72, C2 => n208_port, ZN => 
                           n36_port);
   U99 : BUF_X1 port map( A => b(4), Z => n225_port);
   U100 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => o(0));
   U101 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => o(7));
   U102 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => o(6));
   U103 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => o(5));
   U104 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => o(4));
   U105 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => o(3));
   U106 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => o(2));
   U107 : NAND2_X1 port map( A1 => n62_port, A2 => n63_port, ZN => o(1));
   U108 : NAND2_X1 port map( A1 => n72_port, A2 => n73, ZN => o(15));
   U109 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => o(14));
   U110 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => o(13));
   U111 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => o(12));
   U112 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => o(11));
   U113 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => o(10));
   U114 : NAND2_X1 port map( A1 => n16_port, A2 => n17_port, ZN => o(9));
   U115 : NAND2_X1 port map( A1 => n24_port, A2 => n25_port, ZN => o(8));
   U116 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => o(31));
   U117 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => o(30));
   U118 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => o(29));
   U119 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => o(28));
   U120 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => o(27));
   U121 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => o(26));
   U122 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => o(25));
   U123 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => o(24));
   U124 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => o(23));
   U125 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => o(22));
   U126 : NAND2_X1 port map( A1 => n58_port, A2 => n59_port, ZN => o(21));
   U127 : NAND2_X1 port map( A1 => n60_port, A2 => n61_port, ZN => o(20));
   U128 : NAND2_X1 port map( A1 => n64_port, A2 => n65_port, ZN => o(19));
   U129 : NAND2_X1 port map( A1 => n66_port, A2 => n67_port, ZN => o(18));
   U130 : NAND2_X1 port map( A1 => n68_port, A2 => n69_port, ZN => o(17));
   U131 : NAND2_X1 port map( A1 => n70_port, A2 => n71_port, ZN => o(16));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity DIVIDER_N_op32 is

   port( CLK, START, RESET : in std_logic;  BUSY : out std_logic;  DIVIDEND, 
         DIVISOR : in std_logic_vector (31 downto 0);  QUOTIENT, RESIDUAL : out
         std_logic_vector (31 downto 0));

end DIVIDER_N_op32;

architecture SYN_asd of DIVIDER_N_op32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DIVIDER_N_op32_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component DIVIDER_N_op32_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal RESI_2_31_port, RESI_2_30_port, RESI_2_29_port, RESI_2_28_port, 
      RESI_2_27_port, RESI_2_26_port, RESI_2_25_port, RESI_2_24_port, 
      RESI_2_23_port, RESI_2_22_port, RESI_2_21_port, RESI_2_20_port, 
      RESI_2_19_port, RESI_2_18_port, RESI_2_17_port, RESI_2_16_port, 
      RESI_2_15_port, RESI_2_14_port, RESI_2_13_port, RESI_2_12_port, 
      RESI_2_11_port, RESI_2_10_port, RESI_2_9_port, RESI_2_8_port, 
      RESI_2_7_port, RESI_2_6_port, RESI_2_5_port, RESI_2_4_port, RESI_2_3_port
      , RESI_2_2_port, RESI_2_1_port, RESI_ES_31_port, RESI_ES_30_port, 
      RESI_ES_29_port, RESI_ES_28_port, RESI_ES_27_port, RESI_ES_26_port, 
      RESI_ES_25_port, RESI_ES_24_port, RESI_ES_23_port, RESI_ES_22_port, 
      RESI_ES_21_port, RESI_ES_20_port, RESI_ES_19_port, RESI_ES_18_port, 
      RESI_ES_17_port, RESI_ES_16_port, RESI_ES_15_port, RESI_ES_14_port, 
      RESI_ES_13_port, RESI_ES_12_port, RESI_ES_11_port, RESI_ES_10_port, 
      RESI_ES_9_port, RESI_ES_8_port, RESI_ES_7_port, RESI_ES_6_port, 
      RESI_ES_5_port, RESI_ES_4_port, RESI_ES_3_port, RESI_ES_2_port, 
      RESI_ES_1_port, RESI_ES_0_port, count_31_port, count_30_port, 
      count_29_port, count_28_port, count_27_port, count_26_port, count_25_port
      , count_24_port, count_23_port, count_22_port, count_21_port, 
      count_20_port, count_19_port, count_18_port, count_17_port, count_16_port
      , count_15_port, count_14_port, count_13_port, count_12_port, 
      count_11_port, count_10_port, count_9_port, count_8_port, count_7_port, 
      count_6_port, count_5_port, count_4_port, count_3_port, count_2_port, 
      count_1_port, count_0_port, flag, N172, N173, N174, N175, N176, N177, 
      N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, 
      N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, 
      N202, N203, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, 
      N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, 
      N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172_port, n173_port, n174_port, n175_port, n176_port, 
      n177_port, n178_port, n179_port, n180_port, n181_port, n182_port, 
      n183_port, n184_port, n185_port, n186_port, n187_port, n188_port, 
      n189_port, n190_port, n191_port, n192_port, n193_port, n194_port, 
      n195_port, n196_port, n197_port, n198_port, n199_port, n200_port, 
      n201_port, n202_port, n203_port, n204, n205, n206, n207, n208, n209, n210
      , n244, n245, n246, n248, n249, n250, n251, n252, n253, n254, n255, n256,
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431_port, n432_port, n433_port, 
      n434_port, n435_port, n436_port, n437_port, n438_port, n439_port, 
      n440_port, n441_port, n442_port, n443_port, n444_port, n445_port, 
      n446_port, n447_port, n448_port, n449_port, n450_port, n451_port, 
      n452_port, n453_port, n454_port, n455_port, n456_port, n457_port, 
      n458_port, n459_port, n460_port, n461_port, n462_port, n463, n464, n465, 
      n466, n467, n468, n471, net88277, net88279, net88280, net88281, net88282,
      net88283, net88284, net88285, net88286, net88287, net88288, net88289, 
      net88290, net88291, net88292, net88293, net88294, net88295, net88296, 
      net88297, net88298, net88299, net88300, net88301, net88302, net88303, 
      net88304, net88305, net88338, net166327, n1, n4, n74, n75, n76, n79, n112
      , n113, n114, n116, n117, n119, n121, n123, n125, n127, n129, n131, n133,
      n135, n137, n139, n141, n211, n213, n215, n217, n219, n221, n223, n225, 
      n227, n229, n231, n233, n235, n237, n239, n241, n247, n469, n470, n472, 
      n473, n474, n475, n476, n477, n478, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, 
      n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054 : std_logic;

begin
   
   flag_reg : DFFS_X1 port map( D => n817, CK => n880, SN => n852, Q => flag, 
                           QN => net88338);
   BUSY_reg : DFFS_X1 port map( D => n818, CK => n880, SN => n853, Q => BUSY, 
                           QN => n468);
   QUOTIENT_inter_reg_0_inst : DFF_X1 port map( D => n463, CK => n882, Q => 
                           n_1023, QN => n775);
   QUOTIENT_inter_reg_1_inst : DFF_X1 port map( D => n462_port, CK => n883, Q 
                           => n_1024, QN => n791);
   QUOTIENT_inter_reg_2_inst : DFF_X1 port map( D => n461_port, CK => n882, Q 
                           => n_1025, QN => n776);
   QUOTIENT_inter_reg_3_inst : DFF_X1 port map( D => n460_port, CK => n882, Q 
                           => n_1026, QN => n792);
   QUOTIENT_inter_reg_4_inst : DFF_X1 port map( D => n459_port, CK => n882, Q 
                           => n_1027, QN => n777);
   QUOTIENT_inter_reg_5_inst : DFF_X1 port map( D => n458_port, CK => n883, Q 
                           => n_1028, QN => n793);
   QUOTIENT_inter_reg_6_inst : DFF_X1 port map( D => n457_port, CK => n882, Q 
                           => n_1029, QN => n778);
   QUOTIENT_inter_reg_7_inst : DFF_X1 port map( D => n456_port, CK => n883, Q 
                           => n_1030, QN => n794);
   QUOTIENT_inter_reg_8_inst : DFF_X1 port map( D => n455_port, CK => n881, Q 
                           => n_1031, QN => n779);
   QUOTIENT_inter_reg_9_inst : DFF_X1 port map( D => n454_port, CK => n883, Q 
                           => n_1032, QN => n795);
   QUOTIENT_inter_reg_10_inst : DFF_X1 port map( D => n453_port, CK => n882, Q 
                           => n_1033, QN => n780);
   QUOTIENT_inter_reg_11_inst : DFF_X1 port map( D => n452_port, CK => n882, Q 
                           => n_1034, QN => n796);
   QUOTIENT_inter_reg_12_inst : DFF_X1 port map( D => n451_port, CK => n882, Q 
                           => n_1035, QN => n781);
   QUOTIENT_inter_reg_13_inst : DFF_X1 port map( D => n450_port, CK => n881, Q 
                           => n_1036, QN => n797);
   QUOTIENT_inter_reg_14_inst : DFF_X1 port map( D => n449_port, CK => n882, Q 
                           => n_1037, QN => n782);
   QUOTIENT_inter_reg_15_inst : DFF_X1 port map( D => n448_port, CK => n883, Q 
                           => n_1038, QN => n798);
   QUOTIENT_inter_reg_16_inst : DFF_X1 port map( D => n447_port, CK => n881, Q 
                           => n_1039, QN => n783);
   QUOTIENT_inter_reg_17_inst : DFF_X1 port map( D => n446_port, CK => n883, Q 
                           => n_1040, QN => n799);
   QUOTIENT_inter_reg_18_inst : DFF_X1 port map( D => n445_port, CK => n881, Q 
                           => n_1041, QN => n784);
   QUOTIENT_inter_reg_19_inst : DFF_X1 port map( D => n444_port, CK => n883, Q 
                           => n_1042, QN => n800);
   QUOTIENT_inter_reg_20_inst : DFF_X1 port map( D => n443_port, CK => n881, Q 
                           => n_1043, QN => n785);
   QUOTIENT_inter_reg_21_inst : DFF_X1 port map( D => n442_port, CK => n883, Q 
                           => n_1044, QN => n801);
   QUOTIENT_inter_reg_22_inst : DFF_X1 port map( D => n441_port, CK => n881, Q 
                           => n_1045, QN => n786);
   QUOTIENT_inter_reg_23_inst : DFF_X1 port map( D => n440_port, CK => n881, Q 
                           => n_1046, QN => n802);
   QUOTIENT_inter_reg_24_inst : DFF_X1 port map( D => n439_port, CK => n881, Q 
                           => n_1047, QN => n787);
   QUOTIENT_inter_reg_25_inst : DFF_X1 port map( D => n438_port, CK => n883, Q 
                           => n_1048, QN => n803);
   QUOTIENT_inter_reg_26_inst : DFF_X1 port map( D => n437_port, CK => n881, Q 
                           => n_1049, QN => n788);
   QUOTIENT_inter_reg_27_inst : DFF_X1 port map( D => n436_port, CK => n881, Q 
                           => n_1050, QN => n804);
   QUOTIENT_inter_reg_28_inst : DFF_X1 port map( D => n435_port, CK => n880, Q 
                           => n_1051, QN => n789);
   QUOTIENT_inter_reg_29_inst : DFF_X1 port map( D => n434_port, CK => n882, Q 
                           => n_1052, QN => n805);
   QUOTIENT_inter_reg_30_inst : DFF_X1 port map( D => n433_port, CK => n881, Q 
                           => n_1053, QN => n790);
   QUOTIENT_inter_reg_31_inst : DFF_X1 port map( D => n432_port, CK => n882, Q 
                           => n_1054, QN => n806);
   QUOTIENT_reg_31_inst : DFFR_X1 port map( D => n431_port, CK => n872, RN => 
                           n854, Q => QUOTIENT(31), QN => n210);
   QUOTIENT_reg_30_inst : DFFR_X1 port map( D => n430, CK => n872, RN => n857, 
                           Q => QUOTIENT(30), QN => n209);
   QUOTIENT_reg_29_inst : DFFR_X1 port map( D => n429, CK => n872, RN => n857, 
                           Q => QUOTIENT(29), QN => n208);
   QUOTIENT_reg_28_inst : DFFR_X1 port map( D => n428, CK => n872, RN => n857, 
                           Q => QUOTIENT(28), QN => n207);
   QUOTIENT_reg_27_inst : DFFR_X1 port map( D => n427, CK => n872, RN => n852, 
                           Q => QUOTIENT(27), QN => n206);
   QUOTIENT_reg_26_inst : DFFR_X1 port map( D => n426, CK => n872, RN => n852, 
                           Q => QUOTIENT(26), QN => n205);
   QUOTIENT_reg_25_inst : DFFR_X1 port map( D => n425, CK => n872, RN => n852, 
                           Q => QUOTIENT(25), QN => n204);
   QUOTIENT_reg_24_inst : DFFR_X1 port map( D => n424, CK => n872, RN => n852, 
                           Q => QUOTIENT(24), QN => n203_port);
   QUOTIENT_reg_23_inst : DFFR_X1 port map( D => n423, CK => n872, RN => n852, 
                           Q => QUOTIENT(23), QN => n202_port);
   QUOTIENT_reg_22_inst : DFFR_X1 port map( D => n422, CK => n872, RN => n852, 
                           Q => QUOTIENT(22), QN => n201_port);
   QUOTIENT_reg_21_inst : DFFR_X1 port map( D => n421, CK => n873, RN => n852, 
                           Q => QUOTIENT(21), QN => n200_port);
   QUOTIENT_reg_20_inst : DFFR_X1 port map( D => n420, CK => n873, RN => n852, 
                           Q => QUOTIENT(20), QN => n199_port);
   QUOTIENT_reg_19_inst : DFFR_X1 port map( D => n419, CK => n873, RN => n852, 
                           Q => QUOTIENT(19), QN => n198_port);
   QUOTIENT_reg_18_inst : DFFR_X1 port map( D => n418, CK => n873, RN => n852, 
                           Q => QUOTIENT(18), QN => n197_port);
   QUOTIENT_reg_17_inst : DFFR_X1 port map( D => n417, CK => n873, RN => n852, 
                           Q => QUOTIENT(17), QN => n196_port);
   QUOTIENT_reg_16_inst : DFFR_X1 port map( D => n416, CK => n872, RN => n852, 
                           Q => QUOTIENT(16), QN => n195_port);
   QUOTIENT_reg_15_inst : DFFR_X1 port map( D => n415, CK => n873, RN => n857, 
                           Q => QUOTIENT(15), QN => n194_port);
   QUOTIENT_reg_14_inst : DFFR_X1 port map( D => n414, CK => n873, RN => n856, 
                           Q => QUOTIENT(14), QN => n193_port);
   QUOTIENT_reg_13_inst : DFFR_X1 port map( D => n413, CK => n873, RN => n856, 
                           Q => QUOTIENT(13), QN => n192_port);
   QUOTIENT_reg_12_inst : DFFR_X1 port map( D => n412, CK => n873, RN => n856, 
                           Q => QUOTIENT(12), QN => n191_port);
   QUOTIENT_reg_11_inst : DFFR_X1 port map( D => n411, CK => n873, RN => n856, 
                           Q => QUOTIENT(11), QN => n190_port);
   QUOTIENT_reg_10_inst : DFFR_X1 port map( D => n410, CK => n874, RN => n856, 
                           Q => QUOTIENT(10), QN => n189_port);
   QUOTIENT_reg_9_inst : DFFR_X1 port map( D => n409, CK => n874, RN => n856, Q
                           => QUOTIENT(9), QN => n188_port);
   QUOTIENT_reg_8_inst : DFFR_X1 port map( D => n408, CK => n873, RN => n856, Q
                           => QUOTIENT(8), QN => n187_port);
   QUOTIENT_reg_7_inst : DFFR_X1 port map( D => n407, CK => n874, RN => n856, Q
                           => QUOTIENT(7), QN => n186_port);
   QUOTIENT_reg_6_inst : DFFR_X1 port map( D => n406, CK => n874, RN => n856, Q
                           => QUOTIENT(6), QN => n185_port);
   QUOTIENT_reg_5_inst : DFFR_X1 port map( D => n405, CK => n874, RN => n856, Q
                           => QUOTIENT(5), QN => n184_port);
   QUOTIENT_reg_4_inst : DFFR_X1 port map( D => n404, CK => n874, RN => n856, Q
                           => QUOTIENT(4), QN => n183_port);
   QUOTIENT_reg_3_inst : DFFR_X1 port map( D => n403, CK => n874, RN => n853, Q
                           => QUOTIENT(3), QN => n182_port);
   QUOTIENT_reg_2_inst : DFFR_X1 port map( D => n402, CK => n874, RN => n853, Q
                           => QUOTIENT(2), QN => n181_port);
   QUOTIENT_reg_1_inst : DFFR_X1 port map( D => n401, CK => n874, RN => n853, Q
                           => QUOTIENT(1), QN => n180_port);
   QUOTIENT_reg_0_inst : DFFR_X1 port map( D => n400, CK => n880, RN => n853, Q
                           => QUOTIENT(0), QN => n179_port);
   RESIDUAL_reg_11_inst : DFFR_X1 port map( D => n351, CK => n879, RN => n853, 
                           Q => RESIDUAL(11), QN => n178_port);
   RESIDUAL_reg_10_inst : DFFR_X1 port map( D => n350, CK => n878, RN => n854, 
                           Q => RESIDUAL(10), QN => n177_port);
   RESIDUAL_reg_9_inst : DFFR_X1 port map( D => n349, CK => n878, RN => n854, Q
                           => RESIDUAL(9), QN => n176_port);
   RESIDUAL_reg_8_inst : DFFR_X1 port map( D => n348, CK => n878, RN => n854, Q
                           => RESIDUAL(8), QN => n175_port);
   RESIDUAL_reg_7_inst : DFFR_X1 port map( D => n347, CK => n878, RN => n854, Q
                           => RESIDUAL(7), QN => n174_port);
   RESIDUAL_reg_6_inst : DFFR_X1 port map( D => n346, CK => n877, RN => n854, Q
                           => RESIDUAL(6), QN => n173_port);
   RESIDUAL_reg_5_inst : DFFR_X1 port map( D => n345, CK => n878, RN => n854, Q
                           => RESIDUAL(5), QN => n172_port);
   RESIDUAL_reg_4_inst : DFFR_X1 port map( D => n344, CK => n878, RN => n854, Q
                           => RESIDUAL(4), QN => n171);
   RESIDUAL_reg_3_inst : DFFR_X1 port map( D => n343, CK => n878, RN => n854, Q
                           => RESIDUAL(3), QN => n170);
   RESIDUAL_reg_2_inst : DFFR_X1 port map( D => n342, CK => n878, RN => n854, Q
                           => RESIDUAL(2), QN => n169);
   RESIDUAL_reg_1_inst : DFFR_X1 port map( D => n341, CK => n878, RN => n854, Q
                           => RESIDUAL(1), QN => n168);
   RESIDUAL_reg_0_inst : DFFR_X1 port map( D => n340, CK => n878, RN => n854, Q
                           => RESIDUAL(0), QN => n167);
   RESIDUAL_reg_12_inst : DFFR_X1 port map( D => n335, CK => n879, RN => n853, 
                           Q => RESIDUAL(12), QN => n166);
   RESIDUAL_reg_13_inst : DFFR_X1 port map( D => n330, CK => n879, RN => n853, 
                           Q => RESIDUAL(13), QN => n165);
   RESIDUAL_reg_14_inst : DFFR_X1 port map( D => n325, CK => n878, RN => n853, 
                           Q => RESIDUAL(14), QN => n164);
   RESIDUAL_reg_15_inst : DFFR_X1 port map( D => n320, CK => n879, RN => n853, 
                           Q => RESIDUAL(15), QN => n163);
   RESIDUAL_reg_16_inst : DFFR_X1 port map( D => n315, CK => n879, RN => n853, 
                           Q => RESIDUAL(16), QN => n162);
   RESIDUAL_reg_17_inst : DFFR_X1 port map( D => n310, CK => n879, RN => n853, 
                           Q => RESIDUAL(17), QN => n161);
   RESIDUAL_reg_18_inst : DFFR_X1 port map( D => n305, CK => n879, RN => n853, 
                           Q => RESIDUAL(18), QN => n160);
   RESIDUAL_reg_19_inst : DFFR_X1 port map( D => n300, CK => n879, RN => n855, 
                           Q => RESIDUAL(19), QN => n159);
   RESIDUAL_reg_20_inst : DFFR_X1 port map( D => n295, CK => n879, RN => n855, 
                           Q => RESIDUAL(20), QN => n158);
   RESIDUAL_reg_21_inst : DFFR_X1 port map( D => n290, CK => n879, RN => n855, 
                           Q => RESIDUAL(21), QN => n157);
   RESIDUAL_reg_22_inst : DFFR_X1 port map( D => n285, CK => n879, RN => n855, 
                           Q => RESIDUAL(22), QN => n156);
   RESIDUAL_reg_23_inst : DFFR_X1 port map( D => n280, CK => n880, RN => n855, 
                           Q => RESIDUAL(23), QN => n155);
   RESIDUAL_reg_24_inst : DFFR_X1 port map( D => n275, CK => n880, RN => n855, 
                           Q => RESIDUAL(24), QN => n154);
   RESIDUAL_reg_25_inst : DFFR_X1 port map( D => n270, CK => n880, RN => n855, 
                           Q => RESIDUAL(25), QN => n153);
   RESIDUAL_reg_26_inst : DFFR_X1 port map( D => n265, CK => n880, RN => n855, 
                           Q => RESIDUAL(26), QN => n152);
   RESIDUAL_reg_27_inst : DFFR_X1 port map( D => n260, CK => n880, RN => n855, 
                           Q => RESIDUAL(27), QN => n151);
   RESIDUAL_reg_28_inst : DFFR_X1 port map( D => n255, CK => n880, RN => n855, 
                           Q => RESIDUAL(28), QN => n150);
   RESIDUAL_reg_29_inst : DFFR_X1 port map( D => n250, CK => n880, RN => n854, 
                           Q => RESIDUAL(29), QN => n149);
   RESIDUAL_reg_30_inst : DFFR_X1 port map( D => n249, CK => n877, RN => n855, 
                           Q => RESIDUAL(30), QN => n148);
   RESIDUAL_reg_31_inst : DFFR_X1 port map( D => n244, CK => n877, RN => n855, 
                           Q => RESIDUAL(31), QN => n147);
   count_reg_0_inst : DFFR_X1 port map( D => N431, CK => n877, RN => n857, Q =>
                           count_0_port, QN => n471);
   count_reg_1_inst : DFFR_X1 port map( D => N432, CK => n874, RN => n853, Q =>
                           count_1_port, QN => n146);
   count_reg_2_inst : DFFR_X1 port map( D => N433, CK => n875, RN => n855, Q =>
                           count_2_port, QN => n145);
   count_reg_3_inst : DFFR_X1 port map( D => N434, CK => n875, RN => n852, Q =>
                           count_3_port, QN => n144);
   count_reg_4_inst : DFFR_X1 port map( D => N435, CK => n875, RN => n857, Q =>
                           count_4_port, QN => n143);
   count_reg_5_inst : DFFR_X1 port map( D => N436, CK => n875, RN => n857, Q =>
                           count_5_port, QN => net88305);
   count_reg_6_inst : DFFR_X1 port map( D => N437, CK => n875, RN => n857, Q =>
                           count_6_port, QN => net88304);
   count_reg_7_inst : DFFR_X1 port map( D => N438, CK => n875, RN => n857, Q =>
                           count_7_port, QN => net88303);
   count_reg_8_inst : DFFR_X1 port map( D => N439, CK => n875, RN => n856, Q =>
                           count_8_port, QN => net88302);
   count_reg_9_inst : DFFR_X1 port map( D => N440, CK => n874, RN => n857, Q =>
                           count_9_port, QN => net88301);
   count_reg_10_inst : DFFR_X1 port map( D => N441, CK => n875, RN => n857, Q 
                           => count_10_port, QN => net88300);
   count_reg_11_inst : DFFR_X1 port map( D => N442, CK => n875, RN => n857, Q 
                           => count_11_port, QN => net88299);
   count_reg_12_inst : DFFR_X1 port map( D => N443, CK => n875, RN => n856, Q 
                           => count_12_port, QN => net88298);
   count_reg_13_inst : DFFR_X1 port map( D => N444, CK => n876, RN => n855, Q 
                           => count_13_port, QN => net88297);
   count_reg_14_inst : DFFR_X1 port map( D => N445, CK => n876, RN => n854, Q 
                           => count_14_port, QN => net88296);
   count_reg_15_inst : DFFR_X1 port map( D => N446, CK => n876, RN => n853, Q 
                           => count_15_port, QN => net88295);
   count_reg_16_inst : DFFR_X1 port map( D => N447, CK => n876, RN => n853, Q 
                           => count_16_port, QN => net88294);
   count_reg_17_inst : DFFR_X1 port map( D => N448, CK => n875, RN => n852, Q 
                           => count_17_port, QN => net88293);
   count_reg_18_inst : DFFR_X1 port map( D => N449, CK => n876, RN => n857, Q 
                           => count_18_port, QN => net88292);
   count_reg_19_inst : DFFR_X1 port map( D => N450, CK => n876, RN => n855, Q 
                           => count_19_port, QN => net88291);
   count_reg_20_inst : DFFR_X1 port map( D => N451, CK => n876, RN => n852, Q 
                           => count_20_port, QN => net88290);
   count_reg_21_inst : DFFR_X1 port map( D => N452, CK => n876, RN => n856, Q 
                           => count_21_port, QN => net88289);
   count_reg_22_inst : DFFR_X1 port map( D => N453, CK => n876, RN => n854, Q 
                           => count_22_port, QN => net88288);
   count_reg_23_inst : DFFR_X1 port map( D => N454, CK => n876, RN => n853, Q 
                           => count_23_port, QN => net88287);
   count_reg_24_inst : DFFR_X1 port map( D => N455, CK => n877, RN => n852, Q 
                           => count_24_port, QN => net88286);
   count_reg_25_inst : DFFR_X1 port map( D => N456, CK => n876, RN => n857, Q 
                           => count_25_port, QN => net88285);
   count_reg_26_inst : DFFR_X1 port map( D => N457, CK => n877, RN => n857, Q 
                           => count_26_port, QN => net88284);
   count_reg_27_inst : DFFR_X1 port map( D => N458, CK => n877, RN => n856, Q 
                           => count_27_port, QN => net88283);
   count_reg_28_inst : DFFR_X1 port map( D => N459, CK => n877, RN => n856, Q 
                           => count_28_port, QN => net88282);
   count_reg_29_inst : DFFR_X1 port map( D => N460, CK => n877, RN => n857, Q 
                           => count_29_port, QN => net88281);
   count_reg_30_inst : DFFR_X1 port map( D => N461, CK => n877, RN => n853, Q 
                           => count_30_port, QN => net88280);
   count_reg_31_inst : DFFR_X1 port map( D => N462, CK => n877, RN => n852, Q 
                           => count_31_port, QN => net88279);
   n1 <= '0';
   n4 <= '0';
   add_61 : DIVIDER_N_op32_DW01_inc_0 port map( A(31) => count_31_port, A(30) 
                           => count_30_port, A(29) => count_29_port, A(28) => 
                           count_28_port, A(27) => count_27_port, A(26) => 
                           count_26_port, A(25) => count_25_port, A(24) => 
                           count_24_port, A(23) => count_23_port, A(22) => 
                           count_22_port, A(21) => count_21_port, A(20) => 
                           count_20_port, A(19) => count_19_port, A(18) => 
                           count_18_port, A(17) => count_17_port, A(16) => 
                           count_16_port, A(15) => count_15_port, A(14) => 
                           count_14_port, A(13) => count_13_port, A(12) => 
                           count_12_port, A(11) => count_11_port, A(10) => 
                           count_10_port, A(9) => count_9_port, A(8) => 
                           count_8_port, A(7) => count_7_port, A(6) => 
                           count_6_port, A(5) => count_5_port, A(4) => 
                           count_4_port, A(3) => count_3_port, A(2) => 
                           count_2_port, A(1) => count_1_port, A(0) => 
                           count_0_port, SUM(31) => N203, SUM(30) => N202, 
                           SUM(29) => N201, SUM(28) => N200, SUM(27) => N199, 
                           SUM(26) => N198, SUM(25) => N197, SUM(24) => N196, 
                           SUM(23) => N195, SUM(22) => N194, SUM(21) => N193, 
                           SUM(20) => N192, SUM(19) => N191, SUM(18) => N190, 
                           SUM(17) => N189, SUM(16) => N188, SUM(15) => N187, 
                           SUM(14) => N186, SUM(13) => N185, SUM(12) => N184, 
                           SUM(11) => N183, SUM(10) => N182, SUM(9) => N181, 
                           SUM(8) => N180, SUM(7) => N179, SUM(6) => N178, 
                           SUM(5) => N177, SUM(4) => N176, SUM(3) => N175, 
                           SUM(2) => N174, SUM(1) => N173, SUM(0) => N172);
   sub_34 : DIVIDER_N_op32_DW01_sub_0 port map( A(31) => RESI_2_31_port, A(30) 
                           => RESI_2_30_port, A(29) => RESI_2_29_port, A(28) =>
                           RESI_2_28_port, A(27) => RESI_2_27_port, A(26) => 
                           RESI_2_26_port, A(25) => RESI_2_25_port, A(24) => 
                           RESI_2_24_port, A(23) => RESI_2_23_port, A(22) => 
                           RESI_2_22_port, A(21) => RESI_2_21_port, A(20) => 
                           RESI_2_20_port, A(19) => RESI_2_19_port, A(18) => 
                           RESI_2_18_port, A(17) => RESI_2_17_port, A(16) => 
                           RESI_2_16_port, A(15) => RESI_2_15_port, A(14) => 
                           RESI_2_14_port, A(13) => RESI_2_13_port, A(12) => 
                           RESI_2_12_port, A(11) => RESI_2_11_port, A(10) => 
                           RESI_2_10_port, A(9) => RESI_2_9_port, A(8) => 
                           RESI_2_8_port, A(7) => RESI_2_7_port, A(6) => 
                           RESI_2_6_port, A(5) => RESI_2_5_port, A(4) => 
                           RESI_2_4_port, A(3) => RESI_2_3_port, A(2) => 
                           RESI_2_2_port, A(1) => RESI_2_1_port, A(0) => n1, 
                           B(31) => DIVISOR(31), B(30) => DIVISOR(30), B(29) =>
                           DIVISOR(29), B(28) => DIVISOR(28), B(27) => 
                           DIVISOR(27), B(26) => DIVISOR(26), B(25) => 
                           DIVISOR(25), B(24) => DIVISOR(24), B(23) => 
                           DIVISOR(23), B(22) => DIVISOR(22), B(21) => 
                           DIVISOR(21), B(20) => DIVISOR(20), B(19) => 
                           DIVISOR(19), B(18) => DIVISOR(18), B(17) => 
                           DIVISOR(17), B(16) => DIVISOR(16), B(15) => 
                           DIVISOR(15), B(14) => DIVISOR(14), B(13) => 
                           DIVISOR(13), B(12) => DIVISOR(12), B(11) => 
                           DIVISOR(11), B(10) => DIVISOR(10), B(9) => 
                           DIVISOR(9), B(8) => DIVISOR(8), B(7) => DIVISOR(7), 
                           B(6) => DIVISOR(6), B(5) => DIVISOR(5), B(4) => 
                           DIVISOR(4), B(3) => DIVISOR(3), B(2) => DIVISOR(2), 
                           B(1) => DIVISOR(1), B(0) => DIVISOR(0), CI => n4, 
                           DIFF(31) => RESI_ES_31_port, DIFF(30) => 
                           RESI_ES_30_port, DIFF(29) => RESI_ES_29_port, 
                           DIFF(28) => RESI_ES_28_port, DIFF(27) => 
                           RESI_ES_27_port, DIFF(26) => RESI_ES_26_port, 
                           DIFF(25) => RESI_ES_25_port, DIFF(24) => 
                           RESI_ES_24_port, DIFF(23) => RESI_ES_23_port, 
                           DIFF(22) => RESI_ES_22_port, DIFF(21) => 
                           RESI_ES_21_port, DIFF(20) => RESI_ES_20_port, 
                           DIFF(19) => RESI_ES_19_port, DIFF(18) => 
                           RESI_ES_18_port, DIFF(17) => RESI_ES_17_port, 
                           DIFF(16) => RESI_ES_16_port, DIFF(15) => 
                           RESI_ES_15_port, DIFF(14) => RESI_ES_14_port, 
                           DIFF(13) => RESI_ES_13_port, DIFF(12) => 
                           RESI_ES_12_port, DIFF(11) => RESI_ES_11_port, 
                           DIFF(10) => RESI_ES_10_port, DIFF(9) => 
                           RESI_ES_9_port, DIFF(8) => RESI_ES_8_port, DIFF(7) 
                           => RESI_ES_7_port, DIFF(6) => RESI_ES_6_port, 
                           DIFF(5) => RESI_ES_5_port, DIFF(4) => RESI_ES_4_port
                           , DIFF(3) => RESI_ES_3_port, DIFF(2) => 
                           RESI_ES_2_port, DIFF(1) => RESI_ES_1_port, DIFF(0) 
                           => RESI_ES_0_port, CO => net166327);
   RESIDUAL_inter_reg_31_inst : DFFRS_X1 port map( D => n248, CK => n886, RN =>
                           n245, SN => n246, Q => net88277, QN => n807);
   RESIDUAL_inter_reg_0_inst : DFFRS_X1 port map( D => n399, CK => n886, RN => 
                           n396, SN => n397, Q => RESI_2_1_port, QN => n398);
   RESIDUAL_inter_reg_3_inst : DFFRS_X1 port map( D => n387, CK => n886, RN => 
                           n384, SN => n385, Q => RESI_2_4_port, QN => n386);
   RESIDUAL_inter_reg_30_inst : DFFRS_X1 port map( D => n467, CK => n886, RN =>
                           n464, SN => n465, Q => RESI_2_31_port, QN => n466);
   RESIDUAL_inter_reg_11_inst : DFFRS_X1 port map( D => n355, CK => n886, RN =>
                           n352, SN => n353, Q => RESI_2_12_port, QN => n354);
   RESIDUAL_inter_reg_13_inst : DFFRS_X1 port map( D => n334, CK => n886, RN =>
                           n331, SN => n332, Q => RESI_2_14_port, QN => n333);
   RESIDUAL_inter_reg_23_inst : DFFRS_X1 port map( D => n284, CK => n883, RN =>
                           n281, SN => n282, Q => RESI_2_24_port, QN => n283);
   RESIDUAL_inter_reg_25_inst : DFFRS_X1 port map( D => n274, CK => n883, RN =>
                           n271, SN => n272, Q => RESI_2_26_port, QN => n273);
   RESIDUAL_inter_reg_1_inst : DFFRS_X1 port map( D => n395, CK => n885, RN => 
                           n392, SN => n393, Q => RESI_2_2_port, QN => n394);
   RESIDUAL_inter_reg_4_inst : DFFRS_X1 port map( D => n383, CK => n885, RN => 
                           n380, SN => n381, Q => RESI_2_5_port, QN => n382);
   RESIDUAL_inter_reg_15_inst : DFFRS_X1 port map( D => n324, CK => n884, RN =>
                           n321, SN => n322, Q => RESI_2_16_port, QN => n323);
   RESIDUAL_inter_reg_26_inst : DFFRS_X1 port map( D => n269, CK => n885, RN =>
                           n266, SN => n267, Q => RESI_2_27_port, QN => n268);
   RESIDUAL_inter_reg_27_inst : DFFRS_X1 port map( D => n264, CK => n885, RN =>
                           n261, SN => n262, Q => RESI_2_28_port, QN => n263);
   RESIDUAL_inter_reg_2_inst : DFFRS_X1 port map( D => n391, CK => n884, RN => 
                           n388, SN => n389, Q => RESI_2_3_port, QN => n390);
   RESIDUAL_inter_reg_28_inst : DFFRS_X1 port map( D => n259, CK => n885, RN =>
                           n256, SN => n257, Q => RESI_2_29_port, QN => n258);
   RESIDUAL_inter_reg_29_inst : DFFRS_X1 port map( D => n254, CK => n884, RN =>
                           n251, SN => n252, Q => RESI_2_30_port, QN => n253);
   RESIDUAL_inter_reg_5_inst : DFFRS_X1 port map( D => n379, CK => n885, RN => 
                           n376, SN => n377, Q => RESI_2_6_port, QN => n378);
   RESIDUAL_inter_reg_6_inst : DFFRS_X1 port map( D => n375, CK => n885, RN => 
                           n372, SN => n373, Q => RESI_2_7_port, QN => n374);
   RESIDUAL_inter_reg_7_inst : DFFRS_X1 port map( D => n371, CK => n885, RN => 
                           n368, SN => n369, Q => RESI_2_8_port, QN => n370);
   RESIDUAL_inter_reg_8_inst : DFFRS_X1 port map( D => n367, CK => n884, RN => 
                           n364, SN => n365, Q => RESI_2_9_port, QN => n366);
   RESIDUAL_inter_reg_9_inst : DFFRS_X1 port map( D => n363, CK => n885, RN => 
                           n360, SN => n361, Q => RESI_2_10_port, QN => n362);
   RESIDUAL_inter_reg_10_inst : DFFRS_X1 port map( D => n359, CK => n884, RN =>
                           n356, SN => n357, Q => RESI_2_11_port, QN => n358);
   RESIDUAL_inter_reg_12_inst : DFFRS_X1 port map( D => n339, CK => n884, RN =>
                           n336, SN => n337, Q => RESI_2_13_port, QN => n338);
   RESIDUAL_inter_reg_14_inst : DFFRS_X1 port map( D => n329, CK => n884, RN =>
                           n326, SN => n327, Q => RESI_2_15_port, QN => n328);
   RESIDUAL_inter_reg_16_inst : DFFRS_X1 port map( D => n319, CK => n885, RN =>
                           n316, SN => n317, Q => RESI_2_17_port, QN => n318);
   RESIDUAL_inter_reg_17_inst : DFFRS_X1 port map( D => n314, CK => n885, RN =>
                           n311, SN => n312, Q => RESI_2_18_port, QN => n313);
   RESIDUAL_inter_reg_18_inst : DFFRS_X1 port map( D => n309, CK => n884, RN =>
                           n306, SN => n307, Q => RESI_2_19_port, QN => n308);
   RESIDUAL_inter_reg_19_inst : DFFRS_X1 port map( D => n304, CK => n884, RN =>
                           n301, SN => n302, Q => RESI_2_20_port, QN => n303);
   RESIDUAL_inter_reg_20_inst : DFFRS_X1 port map( D => n299, CK => n884, RN =>
                           n296, SN => n297, Q => RESI_2_21_port, QN => n298);
   RESIDUAL_inter_reg_21_inst : DFFRS_X1 port map( D => n294, CK => n884, RN =>
                           n291, SN => n292, Q => RESI_2_22_port, QN => n293);
   RESIDUAL_inter_reg_22_inst : DFFRS_X1 port map( D => n289, CK => n885, RN =>
                           n286, SN => n287, Q => RESI_2_23_port, QN => n288);
   RESIDUAL_inter_reg_24_inst : DFFRS_X1 port map( D => n279, CK => n884, RN =>
                           n276, SN => n277, Q => RESI_2_25_port, QN => n278);
   U3 : INV_X1 port map( A => n842, ZN => n833);
   U4 : BUF_X1 port map( A => n842, Z => n834);
   U7 : BUF_X1 port map( A => n843, Z => n841);
   U8 : BUF_X1 port map( A => n843, Z => n840);
   U9 : BUF_X1 port map( A => n843, Z => n839);
   U10 : BUF_X1 port map( A => n842, Z => n838);
   U11 : BUF_X1 port map( A => n840, Z => n837);
   U12 : BUF_X1 port map( A => n843, Z => n836);
   U13 : BUF_X1 port map( A => n843, Z => n835);
   U14 : BUF_X1 port map( A => n843, Z => n842);
   U15 : INV_X1 port map( A => n832, ZN => n843);
   U16 : INV_X1 port map( A => n829, ZN => n815);
   U17 : INV_X1 port map( A => n830, ZN => n816);
   U18 : BUF_X1 port map( A => n76, Z => n845);
   U19 : BUF_X1 port map( A => n76, Z => n844);
   U20 : BUF_X1 port map( A => n76, Z => n846);
   U21 : BUF_X1 port map( A => n79, Z => n832);
   U22 : NOR2_X1 port map( A1 => n814, A2 => n866, ZN => n79);
   U23 : BUF_X1 port map( A => n75, Z => n847);
   U24 : BUF_X1 port map( A => n75, Z => n848);
   U25 : BUF_X1 port map( A => n113, Z => n812);
   U26 : BUF_X1 port map( A => n113, Z => n811);
   U27 : BUF_X1 port map( A => n113, Z => n810);
   U28 : BUF_X1 port map( A => n113, Z => n809);
   U29 : BUF_X1 port map( A => n113, Z => n808);
   U30 : BUF_X1 port map( A => n75, Z => n849);
   U31 : BUF_X1 port map( A => n831, Z => n829);
   U32 : BUF_X1 port map( A => n831, Z => n824);
   U33 : BUF_X1 port map( A => n851, Z => n866);
   U34 : BUF_X1 port map( A => n830, Z => n817);
   U35 : BUF_X1 port map( A => n824, Z => n818);
   U36 : BUF_X1 port map( A => n850, Z => n862);
   U37 : BUF_X1 port map( A => n850, Z => n860);
   U38 : BUF_X1 port map( A => n851, Z => n863);
   U39 : BUF_X1 port map( A => n851, Z => n864);
   U40 : BUF_X1 port map( A => n850, Z => n861);
   U41 : BUF_X1 port map( A => n850, Z => n859);
   U42 : BUF_X1 port map( A => n850, Z => n858);
   U43 : BUF_X1 port map( A => n851, Z => n865);
   U44 : BUF_X1 port map( A => n831, Z => n826);
   U45 : BUF_X1 port map( A => n831, Z => n827);
   U46 : BUF_X1 port map( A => n831, Z => n825);
   U47 : BUF_X1 port map( A => n831, Z => n828);
   U48 : BUF_X1 port map( A => n851, Z => n867);
   U49 : BUF_X1 port map( A => n830, Z => n822);
   U50 : BUF_X1 port map( A => n830, Z => n819);
   U51 : BUF_X1 port map( A => n830, Z => n823);
   U52 : BUF_X1 port map( A => n830, Z => n820);
   U53 : BUF_X1 port map( A => n828, Z => n821);
   U54 : BUF_X1 port map( A => n831, Z => n830);
   U55 : INV_X1 port map( A => n241, ZN => n76);
   U56 : NOR2_X1 port map( A1 => n112, A2 => RESI_ES_31_port, ZN => n75);
   U57 : NAND2_X1 port map( A1 => n868, A2 => n814, ZN => n113);
   U58 : OAI22_X1 port map( A1 => n835, A2 => n778, B1 => n79, B2 => n794, ZN 
                           => n456_port);
   U59 : OAI22_X1 port map( A1 => n835, A2 => n793, B1 => n832, B2 => n778, ZN 
                           => n457_port);
   U60 : OAI22_X1 port map( A1 => n835, A2 => n777, B1 => n79, B2 => n793, ZN 
                           => n458_port);
   U61 : OAI22_X1 port map( A1 => n835, A2 => n792, B1 => n832, B2 => n777, ZN 
                           => n459_port);
   U62 : OAI22_X1 port map( A1 => n834, A2 => n776, B1 => n79, B2 => n792, ZN 
                           => n460_port);
   U63 : OAI22_X1 port map( A1 => n834, A2 => n791, B1 => n832, B2 => n776, ZN 
                           => n461_port);
   U64 : OAI22_X1 port map( A1 => n775, A2 => n834, B1 => n79, B2 => n791, ZN 
                           => n462_port);
   U65 : OAI22_X1 port map( A1 => RESI_ES_31_port, A2 => n834, B1 => n832, B2 
                           => n775, ZN => n463);
   U66 : OAI22_X1 port map( A1 => n841, A2 => n790, B1 => n833, B2 => n806, ZN 
                           => n432_port);
   U67 : OAI22_X1 port map( A1 => n841, A2 => n805, B1 => n833, B2 => n790, ZN 
                           => n433_port);
   U68 : OAI22_X1 port map( A1 => n841, A2 => n789, B1 => n833, B2 => n805, ZN 
                           => n434_port);
   U69 : OAI22_X1 port map( A1 => n841, A2 => n804, B1 => n833, B2 => n789, ZN 
                           => n435_port);
   U70 : OAI22_X1 port map( A1 => n840, A2 => n788, B1 => n833, B2 => n804, ZN 
                           => n436_port);
   U71 : OAI22_X1 port map( A1 => n840, A2 => n803, B1 => n833, B2 => n788, ZN 
                           => n437_port);
   U72 : OAI22_X1 port map( A1 => n840, A2 => n787, B1 => n833, B2 => n803, ZN 
                           => n438_port);
   U73 : OAI22_X1 port map( A1 => n840, A2 => n802, B1 => n833, B2 => n787, ZN 
                           => n439_port);
   U74 : OAI22_X1 port map( A1 => n839, A2 => n786, B1 => n833, B2 => n802, ZN 
                           => n440_port);
   U75 : OAI22_X1 port map( A1 => n839, A2 => n801, B1 => n833, B2 => n786, ZN 
                           => n441_port);
   U76 : OAI22_X1 port map( A1 => n839, A2 => n785, B1 => n833, B2 => n801, ZN 
                           => n442_port);
   U77 : OAI22_X1 port map( A1 => n839, A2 => n800, B1 => n833, B2 => n785, ZN 
                           => n443_port);
   U78 : OAI22_X1 port map( A1 => n838, A2 => n784, B1 => n79, B2 => n800, ZN 
                           => n444_port);
   U79 : OAI22_X1 port map( A1 => n838, A2 => n799, B1 => n832, B2 => n784, ZN 
                           => n445_port);
   U80 : OAI22_X1 port map( A1 => n838, A2 => n783, B1 => n79, B2 => n799, ZN 
                           => n446_port);
   U81 : OAI22_X1 port map( A1 => n838, A2 => n798, B1 => n832, B2 => n783, ZN 
                           => n447_port);
   U82 : OAI22_X1 port map( A1 => n837, A2 => n782, B1 => n79, B2 => n798, ZN 
                           => n448_port);
   U83 : OAI22_X1 port map( A1 => n837, A2 => n797, B1 => n832, B2 => n782, ZN 
                           => n449_port);
   U84 : OAI22_X1 port map( A1 => n837, A2 => n781, B1 => n79, B2 => n797, ZN 
                           => n450_port);
   U85 : OAI22_X1 port map( A1 => n837, A2 => n796, B1 => n832, B2 => n781, ZN 
                           => n451_port);
   U86 : OAI22_X1 port map( A1 => n836, A2 => n780, B1 => n79, B2 => n796, ZN 
                           => n452_port);
   U87 : OAI22_X1 port map( A1 => n836, A2 => n795, B1 => n832, B2 => n780, ZN 
                           => n453_port);
   U88 : OAI22_X1 port map( A1 => n836, A2 => n779, B1 => n79, B2 => n795, ZN 
                           => n454_port);
   U89 : OAI22_X1 port map( A1 => n836, A2 => n794, B1 => n832, B2 => n779, ZN 
                           => n455_port);
   U90 : NAND2_X1 port map( A1 => RESI_ES_31_port, A2 => n817, ZN => n241);
   U91 : BUF_X1 port map( A => START, Z => n851);
   U92 : BUF_X1 port map( A => START, Z => n850);
   U93 : INV_X1 port map( A => n814, ZN => n831);
   U94 : AND2_X1 port map( A1 => N176, A2 => n828, ZN => N435);
   U95 : AND2_X1 port map( A1 => N175, A2 => n828, ZN => N434);
   U96 : AND2_X1 port map( A1 => N174, A2 => n829, ZN => N433);
   U97 : AND2_X1 port map( A1 => N173, A2 => n829, ZN => N432);
   U98 : AND2_X1 port map( A1 => N202, A2 => n824, ZN => N461);
   U99 : AND2_X1 port map( A1 => N201, A2 => n825, ZN => N460);
   U100 : AND2_X1 port map( A1 => N200, A2 => n825, ZN => N459);
   U101 : AND2_X1 port map( A1 => N199, A2 => n825, ZN => N458);
   U102 : AND2_X1 port map( A1 => N198, A2 => n825, ZN => N457);
   U103 : AND2_X1 port map( A1 => N197, A2 => n825, ZN => N456);
   U104 : AND2_X1 port map( A1 => N196, A2 => n826, ZN => N455);
   U105 : AND2_X1 port map( A1 => N195, A2 => n826, ZN => N454);
   U106 : AND2_X1 port map( A1 => N194, A2 => n826, ZN => N453);
   U107 : AND2_X1 port map( A1 => N193, A2 => n826, ZN => N452);
   U108 : AND2_X1 port map( A1 => N192, A2 => n826, ZN => N451);
   U109 : AND2_X1 port map( A1 => N191, A2 => n826, ZN => N450);
   U110 : AND2_X1 port map( A1 => N190, A2 => n826, ZN => N449);
   U111 : AND2_X1 port map( A1 => N189, A2 => n827, ZN => N448);
   U112 : AND2_X1 port map( A1 => N188, A2 => n827, ZN => N447);
   U113 : AND2_X1 port map( A1 => N187, A2 => n827, ZN => N446);
   U114 : AND2_X1 port map( A1 => N186, A2 => n827, ZN => N445);
   U115 : AND2_X1 port map( A1 => N185, A2 => n827, ZN => N444);
   U116 : AND2_X1 port map( A1 => N184, A2 => n827, ZN => N443);
   U117 : AND2_X1 port map( A1 => N183, A2 => n827, ZN => N442);
   U118 : AND2_X1 port map( A1 => N182, A2 => n825, ZN => N441);
   U119 : AND2_X1 port map( A1 => N181, A2 => n828, ZN => N440);
   U120 : AND2_X1 port map( A1 => N180, A2 => n828, ZN => N439);
   U121 : AND2_X1 port map( A1 => N179, A2 => n828, ZN => N438);
   U122 : AND2_X1 port map( A1 => N178, A2 => n828, ZN => N437);
   U123 : AND2_X1 port map( A1 => N177, A2 => n828, ZN => N436);
   U124 : NOR4_X1 port map( A1 => count_20_port, A2 => count_19_port, A3 => 
                           count_18_port, A4 => count_17_port, ZN => n474);
   U125 : NOR4_X1 port map( A1 => n471, A2 => n146, A3 => n145, A4 => n144, ZN 
                           => n478);
   U126 : NOR4_X1 port map( A1 => count_16_port, A2 => count_15_port, A3 => 
                           count_14_port, A4 => count_13_port, ZN => n473);
   U127 : NOR4_X1 port map( A1 => n143, A2 => count_31_port, A3 => 
                           count_30_port, A4 => count_29_port, ZN => n477);
   U128 : NOR4_X1 port map( A1 => count_12_port, A2 => count_11_port, A3 => 
                           count_10_port, A4 => count_9_port, ZN => n472);
   U129 : NOR4_X1 port map( A1 => count_28_port, A2 => count_27_port, A3 => 
                           count_26_port, A4 => count_25_port, ZN => n476);
   U130 : NOR4_X1 port map( A1 => count_8_port, A2 => count_7_port, A3 => 
                           count_6_port, A4 => count_5_port, ZN => n470);
   U131 : NOR4_X1 port map( A1 => count_24_port, A2 => count_23_port, A3 => 
                           count_22_port, A4 => count_21_port, ZN => n475);
   U132 : OAI22_X1 port map( A1 => n147, A2 => n814, B1 => n813, B2 => n807, ZN
                           => n244);
   U133 : OAI22_X1 port map( A1 => n148, A2 => n112, B1 => n466, B2 => n813, ZN
                           => n249);
   U134 : OAI22_X1 port map( A1 => n149, A2 => n814, B1 => n253, B2 => n813, ZN
                           => n250);
   U135 : OAI22_X1 port map( A1 => n150, A2 => n814, B1 => n258, B2 => n813, ZN
                           => n255);
   U136 : OAI22_X1 port map( A1 => n824, A2 => n807, B1 => n466, B2 => n241, ZN
                           => n248);
   U137 : OAI22_X1 port map( A1 => n210, A2 => n815, B1 => n806, B2 => n808, ZN
                           => n431_port);
   U138 : OAI22_X1 port map( A1 => n179_port, A2 => n816, B1 => n775, B2 => 
                           n810, ZN => n400);
   U139 : OAI22_X1 port map( A1 => n180_port, A2 => n814, B1 => n791, B2 => 
                           n810, ZN => n401);
   U140 : OAI22_X1 port map( A1 => n181_port, A2 => n814, B1 => n776, B2 => 
                           n810, ZN => n402);
   U141 : OAI22_X1 port map( A1 => n182_port, A2 => n815, B1 => n792, B2 => 
                           n810, ZN => n403);
   U142 : OAI22_X1 port map( A1 => n183_port, A2 => n816, B1 => n777, B2 => 
                           n810, ZN => n404);
   U143 : OAI22_X1 port map( A1 => n184_port, A2 => n814, B1 => n793, B2 => 
                           n810, ZN => n405);
   U144 : OAI22_X1 port map( A1 => n185_port, A2 => n815, B1 => n778, B2 => 
                           n810, ZN => n406);
   U145 : OAI22_X1 port map( A1 => n186_port, A2 => n815, B1 => n794, B2 => 
                           n810, ZN => n407);
   U146 : OAI22_X1 port map( A1 => n187_port, A2 => n816, B1 => n779, B2 => 
                           n809, ZN => n408);
   U147 : OAI22_X1 port map( A1 => n188_port, A2 => n815, B1 => n795, B2 => 
                           n809, ZN => n409);
   U148 : OAI22_X1 port map( A1 => n189_port, A2 => n815, B1 => n780, B2 => 
                           n809, ZN => n410);
   U149 : OAI22_X1 port map( A1 => n190_port, A2 => n815, B1 => n796, B2 => 
                           n809, ZN => n411);
   U150 : OAI22_X1 port map( A1 => n191_port, A2 => n815, B1 => n781, B2 => 
                           n809, ZN => n412);
   U151 : OAI22_X1 port map( A1 => n192_port, A2 => n815, B1 => n797, B2 => 
                           n809, ZN => n413);
   U152 : OAI22_X1 port map( A1 => n193_port, A2 => n815, B1 => n782, B2 => 
                           n809, ZN => n414);
   U153 : OAI22_X1 port map( A1 => n194_port, A2 => n815, B1 => n798, B2 => 
                           n809, ZN => n415);
   U154 : OAI22_X1 port map( A1 => n195_port, A2 => n814, B1 => n783, B2 => 
                           n809, ZN => n416);
   U155 : OAI22_X1 port map( A1 => n196_port, A2 => n815, B1 => n799, B2 => 
                           n809, ZN => n417);
   U156 : OAI22_X1 port map( A1 => n197_port, A2 => n815, B1 => n784, B2 => 
                           n809, ZN => n418);
   U157 : OAI22_X1 port map( A1 => n198_port, A2 => n815, B1 => n800, B2 => 
                           n809, ZN => n419);
   U158 : OAI22_X1 port map( A1 => n199_port, A2 => n815, B1 => n785, B2 => 
                           n808, ZN => n420);
   U159 : OAI22_X1 port map( A1 => n200_port, A2 => n815, B1 => n801, B2 => 
                           n808, ZN => n421);
   U160 : OAI22_X1 port map( A1 => n201_port, A2 => n816, B1 => n786, B2 => 
                           n808, ZN => n422);
   U161 : OAI22_X1 port map( A1 => n202_port, A2 => n815, B1 => n802, B2 => 
                           n808, ZN => n423);
   U162 : OAI22_X1 port map( A1 => n203_port, A2 => n815, B1 => n787, B2 => 
                           n808, ZN => n424);
   U163 : OAI22_X1 port map( A1 => n204, A2 => n816, B1 => n803, B2 => n808, ZN
                           => n425);
   U164 : OAI22_X1 port map( A1 => n205, A2 => n814, B1 => n788, B2 => n808, ZN
                           => n426);
   U165 : OAI22_X1 port map( A1 => n206, A2 => n814, B1 => n804, B2 => n808, ZN
                           => n427);
   U166 : OAI22_X1 port map( A1 => n207, A2 => n816, B1 => n789, B2 => n808, ZN
                           => n428);
   U167 : OAI22_X1 port map( A1 => n208, A2 => n816, B1 => n805, B2 => n808, ZN
                           => n429);
   U168 : OAI22_X1 port map( A1 => n209, A2 => n816, B1 => n790, B2 => n808, ZN
                           => n430);
   U169 : OAI22_X1 port map( A1 => n167, A2 => n112, B1 => n398, B2 => n811, ZN
                           => n340);
   U170 : OAI22_X1 port map( A1 => n151, A2 => n112, B1 => n263, B2 => n812, ZN
                           => n260);
   U171 : OAI22_X1 port map( A1 => n152, A2 => n112, B1 => n268, B2 => n812, ZN
                           => n265);
   U172 : OAI22_X1 port map( A1 => n153, A2 => n816, B1 => n273, B2 => n812, ZN
                           => n270);
   U173 : OAI22_X1 port map( A1 => n154, A2 => n816, B1 => n278, B2 => n812, ZN
                           => n275);
   U174 : OAI22_X1 port map( A1 => n155, A2 => n816, B1 => n283, B2 => n812, ZN
                           => n280);
   U175 : OAI22_X1 port map( A1 => n156, A2 => n816, B1 => n288, B2 => n812, ZN
                           => n285);
   U176 : OAI22_X1 port map( A1 => n157, A2 => n816, B1 => n293, B2 => n812, ZN
                           => n290);
   U177 : OAI22_X1 port map( A1 => n158, A2 => n816, B1 => n298, B2 => n812, ZN
                           => n295);
   U178 : OAI22_X1 port map( A1 => n159, A2 => n816, B1 => n303, B2 => n812, ZN
                           => n300);
   U179 : OAI22_X1 port map( A1 => n160, A2 => n816, B1 => n308, B2 => n812, ZN
                           => n305);
   U180 : OAI22_X1 port map( A1 => n161, A2 => n816, B1 => n313, B2 => n812, ZN
                           => n310);
   U181 : OAI22_X1 port map( A1 => n162, A2 => n816, B1 => n318, B2 => n812, ZN
                           => n315);
   U182 : OAI22_X1 port map( A1 => n163, A2 => n816, B1 => n323, B2 => n811, ZN
                           => n320);
   U183 : OAI22_X1 port map( A1 => n164, A2 => n816, B1 => n328, B2 => n811, ZN
                           => n325);
   U184 : OAI22_X1 port map( A1 => n165, A2 => n814, B1 => n333, B2 => n811, ZN
                           => n330);
   U185 : OAI22_X1 port map( A1 => n166, A2 => n112, B1 => n338, B2 => n811, ZN
                           => n335);
   U186 : OAI22_X1 port map( A1 => n168, A2 => n814, B1 => n394, B2 => n811, ZN
                           => n341);
   U187 : OAI22_X1 port map( A1 => n169, A2 => n112, B1 => n390, B2 => n811, ZN
                           => n342);
   U188 : OAI22_X1 port map( A1 => n170, A2 => n814, B1 => n386, B2 => n811, ZN
                           => n343);
   U189 : OAI22_X1 port map( A1 => n171, A2 => n112, B1 => n382, B2 => n811, ZN
                           => n344);
   U190 : OAI22_X1 port map( A1 => n172_port, A2 => n814, B1 => n378, B2 => 
                           n811, ZN => n345);
   U191 : OAI22_X1 port map( A1 => n173_port, A2 => n112, B1 => n374, B2 => 
                           n811, ZN => n346);
   U192 : OAI22_X1 port map( A1 => n174_port, A2 => n814, B1 => n370, B2 => 
                           n811, ZN => n347);
   U193 : OAI22_X1 port map( A1 => n175_port, A2 => n112, B1 => n366, B2 => 
                           n810, ZN => n348);
   U194 : OAI22_X1 port map( A1 => n176_port, A2 => n814, B1 => n362, B2 => 
                           n810, ZN => n349);
   U195 : OAI22_X1 port map( A1 => n177_port, A2 => n112, B1 => n358, B2 => 
                           n810, ZN => n350);
   U196 : OAI22_X1 port map( A1 => n178_port, A2 => n815, B1 => n354, B2 => 
                           n810, ZN => n351);
   U197 : OAI21_X1 port map( B1 => n273, B2 => n823, A => n231, ZN => n274);
   U198 : AOI22_X1 port map( A1 => RESI_ES_25_port, A2 => n847, B1 => n846, B2 
                           => RESI_2_25_port, ZN => n231);
   U199 : OAI21_X1 port map( B1 => n278, B2 => n822, A => n229, ZN => n279);
   U200 : AOI22_X1 port map( A1 => RESI_ES_24_port, A2 => n847, B1 => n846, B2 
                           => RESI_2_24_port, ZN => n229);
   U201 : OAI21_X1 port map( B1 => n283, B2 => n824, A => n227, ZN => n284);
   U202 : AOI22_X1 port map( A1 => RESI_ES_23_port, A2 => n847, B1 => n845, B2 
                           => RESI_2_23_port, ZN => n227);
   U203 : OAI21_X1 port map( B1 => n288, B2 => n822, A => n225, ZN => n289);
   U204 : AOI22_X1 port map( A1 => RESI_ES_22_port, A2 => n847, B1 => n845, B2 
                           => RESI_2_22_port, ZN => n225);
   U205 : OAI21_X1 port map( B1 => n293, B2 => n822, A => n223, ZN => n294);
   U206 : AOI22_X1 port map( A1 => RESI_ES_21_port, A2 => n847, B1 => n845, B2 
                           => RESI_2_21_port, ZN => n223);
   U207 : OAI21_X1 port map( B1 => n298, B2 => n822, A => n221, ZN => n299);
   U208 : AOI22_X1 port map( A1 => RESI_ES_20_port, A2 => n847, B1 => n845, B2 
                           => RESI_2_20_port, ZN => n221);
   U209 : OAI21_X1 port map( B1 => n303, B2 => n821, A => n219, ZN => n304);
   U210 : AOI22_X1 port map( A1 => RESI_ES_19_port, A2 => n847, B1 => n845, B2 
                           => RESI_2_19_port, ZN => n219);
   U211 : OAI21_X1 port map( B1 => n308, B2 => n821, A => n217, ZN => n309);
   U212 : AOI22_X1 port map( A1 => RESI_ES_18_port, A2 => n847, B1 => n845, B2 
                           => RESI_2_18_port, ZN => n217);
   U213 : OAI21_X1 port map( B1 => n313, B2 => n821, A => n215, ZN => n314);
   U214 : AOI22_X1 port map( A1 => RESI_ES_17_port, A2 => n848, B1 => n845, B2 
                           => RESI_2_17_port, ZN => n215);
   U215 : OAI21_X1 port map( B1 => n318, B2 => n824, A => n213, ZN => n319);
   U216 : AOI22_X1 port map( A1 => RESI_ES_16_port, A2 => n848, B1 => n845, B2 
                           => RESI_2_16_port, ZN => n213);
   U217 : OAI21_X1 port map( B1 => n328, B2 => n820, A => n141, ZN => n329);
   U218 : AOI22_X1 port map( A1 => RESI_ES_14_port, A2 => n848, B1 => n845, B2 
                           => RESI_2_14_port, ZN => n141);
   U219 : OAI21_X1 port map( B1 => n333, B2 => n820, A => n139, ZN => n334);
   U220 : AOI22_X1 port map( A1 => RESI_ES_13_port, A2 => n848, B1 => n845, B2 
                           => RESI_2_13_port, ZN => n139);
   U221 : OAI21_X1 port map( B1 => n338, B2 => n820, A => n137, ZN => n339);
   U222 : AOI22_X1 port map( A1 => RESI_ES_12_port, A2 => n848, B1 => n845, B2 
                           => RESI_2_12_port, ZN => n137);
   U223 : OAI21_X1 port map( B1 => n354, B2 => n819, A => n135, ZN => n355);
   U224 : AOI22_X1 port map( A1 => RESI_ES_11_port, A2 => n848, B1 => n844, B2 
                           => RESI_2_11_port, ZN => n135);
   U225 : OAI21_X1 port map( B1 => n358, B2 => n819, A => n133, ZN => n359);
   U226 : AOI22_X1 port map( A1 => RESI_ES_10_port, A2 => n848, B1 => n844, B2 
                           => RESI_2_10_port, ZN => n133);
   U227 : OAI21_X1 port map( B1 => n362, B2 => n819, A => n131, ZN => n363);
   U228 : AOI22_X1 port map( A1 => RESI_ES_9_port, A2 => n848, B1 => n844, B2 
                           => RESI_2_9_port, ZN => n131);
   U229 : OAI21_X1 port map( B1 => n366, B2 => n819, A => n129, ZN => n367);
   U230 : AOI22_X1 port map( A1 => RESI_ES_8_port, A2 => n848, B1 => n844, B2 
                           => RESI_2_8_port, ZN => n129);
   U231 : OAI21_X1 port map( B1 => n370, B2 => n818, A => n127, ZN => n371);
   U232 : AOI22_X1 port map( A1 => RESI_ES_7_port, A2 => n848, B1 => n844, B2 
                           => RESI_2_7_port, ZN => n127);
   U233 : OAI21_X1 port map( B1 => n374, B2 => n818, A => n125, ZN => n375);
   U234 : AOI22_X1 port map( A1 => RESI_ES_6_port, A2 => n848, B1 => n844, B2 
                           => RESI_2_6_port, ZN => n125);
   U235 : OAI21_X1 port map( B1 => n378, B2 => n818, A => n123, ZN => n379);
   U236 : AOI22_X1 port map( A1 => RESI_ES_5_port, A2 => n849, B1 => n844, B2 
                           => RESI_2_5_port, ZN => n123);
   U237 : OAI21_X1 port map( B1 => n253, B2 => n824, A => n239, ZN => n254);
   U238 : AOI22_X1 port map( A1 => RESI_ES_29_port, A2 => n847, B1 => n846, B2 
                           => RESI_2_29_port, ZN => n239);
   U239 : OAI21_X1 port map( B1 => n258, B2 => n823, A => n237, ZN => n259);
   U240 : AOI22_X1 port map( A1 => RESI_ES_28_port, A2 => n847, B1 => n846, B2 
                           => RESI_2_28_port, ZN => n237);
   U241 : OAI21_X1 port map( B1 => n390, B2 => n817, A => n117, ZN => n391);
   U242 : AOI22_X1 port map( A1 => RESI_ES_2_port, A2 => n849, B1 => n844, B2 
                           => RESI_2_2_port, ZN => n117);
   U243 : OAI21_X1 port map( B1 => n263, B2 => n823, A => n235, ZN => n264);
   U244 : AOI22_X1 port map( A1 => RESI_ES_27_port, A2 => n847, B1 => n846, B2 
                           => RESI_2_27_port, ZN => n235);
   U245 : OAI21_X1 port map( B1 => n268, B2 => n823, A => n233, ZN => n269);
   U246 : AOI22_X1 port map( A1 => RESI_ES_26_port, A2 => n847, B1 => n846, B2 
                           => RESI_2_26_port, ZN => n233);
   U247 : OAI21_X1 port map( B1 => n323, B2 => n820, A => n211, ZN => n324);
   U248 : AOI22_X1 port map( A1 => RESI_ES_15_port, A2 => n848, B1 => n845, B2 
                           => RESI_2_15_port, ZN => n211);
   U249 : OAI21_X1 port map( B1 => n382, B2 => n818, A => n121, ZN => n383);
   U250 : AOI22_X1 port map( A1 => RESI_ES_4_port, A2 => n849, B1 => n844, B2 
                           => RESI_2_4_port, ZN => n121);
   U251 : OAI21_X1 port map( B1 => n386, B2 => n821, A => n119, ZN => n387);
   U252 : AOI22_X1 port map( A1 => RESI_ES_3_port, A2 => n849, B1 => n844, B2 
                           => RESI_2_3_port, ZN => n119);
   U253 : OAI21_X1 port map( B1 => n394, B2 => n817, A => n116, ZN => n395);
   U254 : AOI22_X1 port map( A1 => RESI_ES_1_port, A2 => n849, B1 => n844, B2 
                           => RESI_2_1_port, ZN => n116);
   U255 : OAI21_X1 port map( B1 => n466, B2 => n817, A => n74, ZN => n467);
   U256 : AOI22_X1 port map( A1 => RESI_ES_30_port, A2 => n849, B1 => n844, B2 
                           => RESI_2_30_port, ZN => n74);
   U257 : BUF_X1 port map( A => n112, Z => n814);
   U258 : OAI211_X1 port map( C1 => n247, C2 => n469, A => n868, B => flag, ZN 
                           => n112);
   U259 : NAND4_X1 port map( A1 => n475, A2 => n476, A3 => n477, A4 => n478, ZN
                           => n247);
   U260 : NAND4_X1 port map( A1 => n470, A2 => n472, A3 => n473, A4 => n474, ZN
                           => n469);
   U261 : BUF_X1 port map( A => CLK, Z => n869);
   U262 : BUF_X1 port map( A => CLK, Z => n870);
   U263 : NAND2_X1 port map( A1 => DIVIDEND(25), A2 => n864, ZN => n272);
   U264 : NAND2_X1 port map( A1 => DIVIDEND(24), A2 => n864, ZN => n277);
   U265 : NAND2_X1 port map( A1 => DIVIDEND(23), A2 => n864, ZN => n282);
   U266 : NAND2_X1 port map( A1 => DIVIDEND(22), A2 => n863, ZN => n287);
   U267 : NAND2_X1 port map( A1 => DIVIDEND(21), A2 => n863, ZN => n292);
   U268 : NAND2_X1 port map( A1 => DIVIDEND(20), A2 => n863, ZN => n297);
   U269 : NAND2_X1 port map( A1 => DIVIDEND(19), A2 => n862, ZN => n302);
   U270 : NAND2_X1 port map( A1 => DIVIDEND(18), A2 => n862, ZN => n307);
   U271 : NAND2_X1 port map( A1 => DIVIDEND(17), A2 => n862, ZN => n312);
   U272 : NAND2_X1 port map( A1 => DIVIDEND(16), A2 => n862, ZN => n317);
   U273 : NAND2_X1 port map( A1 => DIVIDEND(14), A2 => n861, ZN => n327);
   U274 : NAND2_X1 port map( A1 => DIVIDEND(13), A2 => n861, ZN => n332);
   U275 : NAND2_X1 port map( A1 => DIVIDEND(12), A2 => n861, ZN => n337);
   U276 : NAND2_X1 port map( A1 => DIVIDEND(11), A2 => n860, ZN => n353);
   U277 : NAND2_X1 port map( A1 => DIVIDEND(10), A2 => n860, ZN => n357);
   U278 : NAND2_X1 port map( A1 => DIVIDEND(9), A2 => n860, ZN => n361);
   U279 : NAND2_X1 port map( A1 => DIVIDEND(8), A2 => n860, ZN => n365);
   U280 : NAND2_X1 port map( A1 => DIVIDEND(7), A2 => n859, ZN => n369);
   U281 : NAND2_X1 port map( A1 => DIVIDEND(6), A2 => n859, ZN => n373);
   U282 : NAND2_X1 port map( A1 => DIVIDEND(5), A2 => n859, ZN => n377);
   U283 : NAND2_X1 port map( A1 => DIVIDEND(29), A2 => n865, ZN => n252);
   U284 : NAND2_X1 port map( A1 => DIVIDEND(28), A2 => n865, ZN => n257);
   U285 : NAND2_X1 port map( A1 => DIVIDEND(2), A2 => n858, ZN => n389);
   U286 : NAND2_X1 port map( A1 => DIVIDEND(30), A2 => n863, ZN => n465);
   U287 : NAND2_X1 port map( A1 => DIVIDEND(27), A2 => n865, ZN => n262);
   U288 : NAND2_X1 port map( A1 => DIVIDEND(26), A2 => n864, ZN => n267);
   U289 : NAND2_X1 port map( A1 => DIVIDEND(15), A2 => n861, ZN => n322);
   U290 : NAND2_X1 port map( A1 => DIVIDEND(4), A2 => n859, ZN => n381);
   U291 : NAND2_X1 port map( A1 => DIVIDEND(3), A2 => n858, ZN => n385);
   U292 : NAND2_X1 port map( A1 => DIVIDEND(1), A2 => n858, ZN => n393);
   U293 : NAND2_X1 port map( A1 => DIVIDEND(0), A2 => n858, ZN => n397);
   U294 : NAND2_X1 port map( A1 => DIVIDEND(31), A2 => n865, ZN => n246);
   U295 : INV_X1 port map( A => n114, ZN => n399);
   U296 : AOI22_X1 port map( A1 => RESI_ES_0_port, A2 => n849, B1 => n814, B2 
                           => RESI_2_1_port, ZN => n114);
   U297 : OR2_X1 port map( A1 => n853, A2 => DIVIDEND(21), ZN => n291);
   U298 : OR2_X1 port map( A1 => n852, A2 => DIVIDEND(20), ZN => n296);
   U299 : OR2_X1 port map( A1 => n855, A2 => DIVIDEND(19), ZN => n301);
   U300 : OR2_X1 port map( A1 => n856, A2 => DIVIDEND(18), ZN => n306);
   U301 : OR2_X1 port map( A1 => n857, A2 => DIVIDEND(17), ZN => n311);
   U302 : OR2_X1 port map( A1 => n853, A2 => DIVIDEND(16), ZN => n316);
   U303 : OR2_X1 port map( A1 => n856, A2 => DIVIDEND(14), ZN => n326);
   U304 : OR2_X1 port map( A1 => n855, A2 => DIVIDEND(13), ZN => n331);
   U305 : OR2_X1 port map( A1 => n854, A2 => DIVIDEND(12), ZN => n336);
   U306 : OR2_X1 port map( A1 => n857, A2 => DIVIDEND(11), ZN => n352);
   U307 : OR2_X1 port map( A1 => n852, A2 => DIVIDEND(10), ZN => n356);
   U308 : OR2_X1 port map( A1 => n855, A2 => DIVIDEND(9), ZN => n360);
   U309 : OR2_X1 port map( A1 => n854, A2 => DIVIDEND(8), ZN => n364);
   U310 : OR2_X1 port map( A1 => n854, A2 => DIVIDEND(7), ZN => n368);
   U311 : OR2_X1 port map( A1 => n857, A2 => DIVIDEND(6), ZN => n372);
   U312 : OR2_X1 port map( A1 => n857, A2 => DIVIDEND(5), ZN => n376);
   U313 : OR2_X1 port map( A1 => n856, A2 => DIVIDEND(2), ZN => n388);
   U314 : OR2_X1 port map( A1 => n855, A2 => DIVIDEND(30), ZN => n464);
   U315 : OR2_X1 port map( A1 => n854, A2 => DIVIDEND(15), ZN => n321);
   U316 : OR2_X1 port map( A1 => n852, A2 => DIVIDEND(4), ZN => n380);
   U317 : OR2_X1 port map( A1 => n854, A2 => DIVIDEND(3), ZN => n384);
   U318 : OR2_X1 port map( A1 => n854, A2 => DIVIDEND(1), ZN => n392);
   U319 : OR2_X1 port map( A1 => n855, A2 => DIVIDEND(0), ZN => n396);
   U320 : OR2_X1 port map( A1 => n857, A2 => DIVIDEND(31), ZN => n245);
   U321 : OR2_X1 port map( A1 => n855, A2 => DIVIDEND(25), ZN => n271);
   U322 : OR2_X1 port map( A1 => n853, A2 => DIVIDEND(24), ZN => n276);
   U323 : OR2_X1 port map( A1 => n857, A2 => DIVIDEND(23), ZN => n281);
   U324 : OR2_X1 port map( A1 => n856, A2 => DIVIDEND(22), ZN => n286);
   U325 : OR2_X1 port map( A1 => n856, A2 => DIVIDEND(29), ZN => n251);
   U326 : OR2_X1 port map( A1 => n854, A2 => DIVIDEND(28), ZN => n256);
   U327 : OR2_X1 port map( A1 => n855, A2 => DIVIDEND(27), ZN => n261);
   U328 : OR2_X1 port map( A1 => n856, A2 => DIVIDEND(26), ZN => n266);
   U329 : BUF_X1 port map( A => CLK, Z => n871);
   U330 : AND2_X1 port map( A1 => N203, A2 => n825, ZN => N462);
   U331 : AND2_X1 port map( A1 => N172, A2 => n829, ZN => N431);
   U332 : CLKBUF_X1 port map( A => n113, Z => n813);
   U333 : INV_X1 port map( A => n866, ZN => n852);
   U334 : INV_X1 port map( A => n866, ZN => n853);
   U335 : INV_X1 port map( A => n866, ZN => n854);
   U336 : INV_X1 port map( A => n866, ZN => n855);
   U337 : INV_X1 port map( A => n866, ZN => n856);
   U338 : INV_X1 port map( A => n867, ZN => n857);
   U339 : INV_X1 port map( A => RESET, ZN => n868);
   U340 : CLKBUF_X1 port map( A => n869, Z => n872);
   U341 : CLKBUF_X1 port map( A => n869, Z => n873);
   U342 : CLKBUF_X1 port map( A => n869, Z => n874);
   U343 : CLKBUF_X1 port map( A => n869, Z => n875);
   U344 : CLKBUF_X1 port map( A => n869, Z => n876);
   U345 : CLKBUF_X1 port map( A => n869, Z => n877);
   U346 : CLKBUF_X1 port map( A => n870, Z => n878);
   U347 : CLKBUF_X1 port map( A => n870, Z => n879);
   U348 : CLKBUF_X1 port map( A => n870, Z => n880);
   U349 : CLKBUF_X1 port map( A => n870, Z => n881);
   U350 : CLKBUF_X1 port map( A => n870, Z => n882);
   U351 : CLKBUF_X1 port map( A => n870, Z => n883);
   U352 : CLKBUF_X1 port map( A => n871, Z => n884);
   U353 : CLKBUF_X1 port map( A => n871, Z => n885);
   U354 : CLKBUF_X1 port map( A => n871, Z => n886);

end SYN_asd;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity forwarding_unit is

   port( EX_MEM_write : in std_logic;  EX_MEM_Rd, ID_EX_Rs, ID_EX_Rt : in 
         std_logic_vector (4 downto 0);  MEM_WB_write : in std_logic;  
         MEM_WB_Rd : in std_logic_vector (4 downto 0);  sel_mux_high, 
         sel_mux_low : out std_logic_vector (1 downto 0));

end forwarding_unit;

architecture SYN_Structural of forwarding_unit is

   component cu_lower_mux
      port( EX_MEM_write, MEM_WB_write : in std_logic;  EX_MEM_Rd, ID_EX_Rt, 
            MEM_WB_Rd : in std_logic_vector (4 downto 0);  sel_lower_mux : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component cu_upper_mux
      port( EX_MEM_write, MEM_WB_write : in std_logic;  MEM_WB_Rd, EX_MEM_Rd, 
            ID_EX_Rs : in std_logic_vector (4 downto 0);  sel_upper_mux : out 
            std_logic_vector (1 downto 0));
   end component;

begin
   
   CU_U_M : cu_upper_mux port map( EX_MEM_write => EX_MEM_write, MEM_WB_write 
                           => MEM_WB_write, MEM_WB_Rd(4) => MEM_WB_Rd(4), 
                           MEM_WB_Rd(3) => MEM_WB_Rd(3), MEM_WB_Rd(2) => 
                           MEM_WB_Rd(2), MEM_WB_Rd(1) => MEM_WB_Rd(1), 
                           MEM_WB_Rd(0) => MEM_WB_Rd(0), EX_MEM_Rd(4) => 
                           EX_MEM_Rd(4), EX_MEM_Rd(3) => EX_MEM_Rd(3), 
                           EX_MEM_Rd(2) => EX_MEM_Rd(2), EX_MEM_Rd(1) => 
                           EX_MEM_Rd(1), EX_MEM_Rd(0) => EX_MEM_Rd(0), 
                           ID_EX_Rs(4) => ID_EX_Rs(4), ID_EX_Rs(3) => 
                           ID_EX_Rs(3), ID_EX_Rs(2) => ID_EX_Rs(2), ID_EX_Rs(1)
                           => ID_EX_Rs(1), ID_EX_Rs(0) => ID_EX_Rs(0), 
                           sel_upper_mux(1) => sel_mux_high(1), 
                           sel_upper_mux(0) => sel_mux_high(0));
   CU_L_M : cu_lower_mux port map( EX_MEM_write => EX_MEM_write, MEM_WB_write 
                           => MEM_WB_write, EX_MEM_Rd(4) => EX_MEM_Rd(4), 
                           EX_MEM_Rd(3) => EX_MEM_Rd(3), EX_MEM_Rd(2) => 
                           EX_MEM_Rd(2), EX_MEM_Rd(1) => EX_MEM_Rd(1), 
                           EX_MEM_Rd(0) => EX_MEM_Rd(0), ID_EX_Rt(4) => 
                           ID_EX_Rt(4), ID_EX_Rt(3) => ID_EX_Rt(3), ID_EX_Rt(2)
                           => ID_EX_Rt(2), ID_EX_Rt(1) => ID_EX_Rt(1), 
                           ID_EX_Rt(0) => ID_EX_Rt(0), MEM_WB_Rd(4) => 
                           MEM_WB_Rd(4), MEM_WB_Rd(3) => MEM_WB_Rd(3), 
                           MEM_WB_Rd(2) => MEM_WB_Rd(2), MEM_WB_Rd(1) => 
                           MEM_WB_Rd(1), MEM_WB_Rd(0) => MEM_WB_Rd(0), 
                           sel_lower_mux(1) => sel_mux_low(1), sel_lower_mux(0)
                           => sel_mux_low(0));

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity mux_2_1_5bit is

   port( a, b : in std_logic_vector (4 downto 0);  sel : in std_logic;  o : out
         std_logic_vector (4 downto 0));

end mux_2_1_5bit;

architecture SYN_Behavioral of mux_2_1_5bit is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n8);
   U2 : INV_X1 port map( A => n12, ZN => o(0));
   U3 : AOI22_X1 port map( A1 => a(0), A2 => sel, B1 => b(0), B2 => n8, ZN => 
                           n12);
   U4 : INV_X1 port map( A => n11, ZN => o(1));
   U5 : AOI22_X1 port map( A1 => a(1), A2 => sel, B1 => b(1), B2 => n8, ZN => 
                           n11);
   U6 : INV_X1 port map( A => n10, ZN => o(2));
   U7 : AOI22_X1 port map( A1 => a(2), A2 => sel, B1 => b(2), B2 => n8, ZN => 
                           n10);
   U8 : INV_X1 port map( A => n9, ZN => o(3));
   U9 : AOI22_X1 port map( A1 => a(3), A2 => sel, B1 => b(3), B2 => n8, ZN => 
                           n9);
   U10 : INV_X1 port map( A => n7, ZN => o(4));
   U11 : AOI22_X1 port map( A1 => sel, A2 => a(4), B1 => b(4), B2 => n8, ZN => 
                           n7);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity cu_exe is

   port( reset : in std_logic;  func : in std_logic_vector (10 downto 0);  
         busy_div : in std_logic;  multi_cycle_operation, enable : out 
         std_logic;  sel_signal_5X1 : out std_logic_vector (2 downto 0);  
         sel_signal_2X1, start_div : out std_logic;  cmd_t2 : out 
         std_logic_vector (3 downto 0);  carry_in, left_right, logic_Arith, 
         shift_rot : out std_logic;  sel_comparator : out std_logic_vector (2 
         downto 0));

end cu_exe;

architecture SYN_Behavioral of cu_exe is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, sel_signal_5X1_1_port, sel_signal_5X1_0_port, 
      cmd_t2_3_port, sel_comparator_2_port, sel_comparator_1_port, 
      sel_comparator_0_port, cmd_t2_1_port, sel_signal_5X1_2_port, 
      sel_signal_2X1_port, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n76 : std_logic;

begin
   multi_cycle_operation <= sel_signal_2X1_port;
   sel_signal_5X1 <= ( sel_signal_5X1_2_port, sel_signal_5X1_1_port, 
      sel_signal_5X1_0_port );
   sel_signal_2X1 <= sel_signal_2X1_port;
   cmd_t2 <= ( cmd_t2_3_port, cmd_t2_1_port, cmd_t2_1_port, X_Logic0_port );
   sel_comparator <= ( sel_comparator_2_port, sel_comparator_1_port, 
      sel_comparator_0_port );
   
   X_Logic0_port <= '0';
   U44 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => n18, ZN => 
                           sel_signal_5X1_0_port);
   U45 : NAND3_X1 port map( A1 => n26, A2 => n76, A3 => func(3), ZN => 
                           sel_comparator_1_port);
   U3 : NOR4_X1 port map( A1 => func(6), A2 => func(5), A3 => func(10), A4 => 
                           n40, ZN => n36);
   U4 : NOR2_X1 port map( A1 => n32, A2 => func(1), ZN => n26);
   U5 : INV_X1 port map( A => n37, ZN => n24);
   U6 : NOR3_X1 port map( A1 => n19, A2 => n20, A3 => n21, ZN => 
                           sel_signal_2X1_port);
   U7 : NAND2_X1 port map( A1 => n31, A2 => n26, ZN => n20);
   U8 : NAND2_X1 port map( A1 => n22, A2 => n19, ZN => sel_comparator_0_port);
   U9 : NAND2_X1 port map( A1 => n22, A2 => n21, ZN => sel_comparator_2_port);
   U10 : NOR3_X1 port map( A1 => n14, A2 => reset, A3 => n15, ZN => shift_rot);
   U11 : NOR2_X1 port map( A1 => n19, A2 => n18, ZN => left_right);
   U12 : OAI21_X1 port map( B1 => n33, B2 => n34, A => n76, ZN => n18);
   U13 : INV_X1 port map( A => n15, ZN => n33);
   U14 : NOR4_X1 port map( A1 => n32, A2 => n21, A3 => n14, A4 => n35, ZN => 
                           n34);
   U15 : NAND2_X1 port map( A1 => sel_comparator_2_port, A2 => 
                           sel_comparator_1_port, ZN => sel_signal_5X1_2_port);
   U16 : INV_X1 port map( A => n17, ZN => cmd_t2_1_port);
   U17 : OR3_X1 port map( A1 => func(9), A2 => func(8), A3 => func(7), ZN => 
                           n40);
   U18 : INV_X1 port map( A => func(4), ZN => n39);
   U19 : NOR3_X1 port map( A1 => n32, A2 => func(2), A3 => n14, ZN => n29);
   U20 : NOR2_X1 port map( A1 => func(3), A2 => reset, ZN => n31);
   U21 : INV_X1 port map( A => func(2), ZN => n21);
   U22 : INV_X1 port map( A => func(0), ZN => n19);
   U23 : INV_X1 port map( A => func(1), ZN => n14);
   U24 : INV_X1 port map( A => reset, ZN => n76);
   U25 : INV_X1 port map( A => n28, ZN => n22);
   U26 : NOR3_X1 port map( A1 => n15, A2 => reset, A3 => func(1), ZN => 
                           logic_Arith);
   U27 : NAND2_X1 port map( A1 => n18, A2 => n30, ZN => sel_signal_5X1_1_port);
   U28 : OR3_X1 port map( A1 => n20, A2 => func(0), A3 => n21, ZN => n30);
   U29 : NAND4_X1 port map( A1 => func(1), A2 => func(2), A3 => n31, A4 => n38,
                           ZN => n17);
   U30 : INV_X1 port map( A => n32, ZN => n38);
   U31 : NOR2_X1 port map( A1 => busy_div, A2 => n13, ZN => start_div);
   U32 : INV_X1 port map( A => sel_signal_2X1_port, ZN => n13);
   U33 : OR4_X1 port map( A1 => sel_signal_5X1_1_port, A2 => 
                           sel_signal_5X1_2_port, A3 => cmd_t2_1_port, A4 => 
                           n23, ZN => enable);
   U34 : OR2_X1 port map( A1 => n24, A2 => n25, ZN => n23);
   U35 : NOR3_X1 port map( A1 => n19, A2 => func(2), A3 => n20, ZN => n25);
   U36 : OAI21_X1 port map( B1 => func(0), B2 => n17, A => n16, ZN => 
                           cmd_t2_3_port);
   U37 : NAND2_X1 port map( A1 => n24, A2 => func(0), ZN => n16);
   U38 : INV_X1 port map( A => func(3), ZN => n35);
   U39 : NOR2_X1 port map( A1 => func(0), A2 => n37, ZN => carry_in);
   U40 : NAND2_X1 port map( A1 => n29, A2 => n31, ZN => n37);
   U41 : NAND4_X1 port map( A1 => func(4), A2 => n36, A3 => n21, A4 => n35, ZN 
                           => n15);
   U42 : OAI211_X1 port map( C1 => n29, C2 => n26, A => n76, B => func(3), ZN 
                           => n28);
   U43 : NAND2_X1 port map( A1 => n36, A2 => n39, ZN => n32);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity fetchUnit is

   port( sel0, en0, clock, reset : in std_logic;  fromInstructionMemory, 
         next_PC : in std_logic_vector (31 downto 0);  PcToInstructionMemory, 
         InstructionToDecode, pcToDecode : out std_logic_vector (31 downto 0));

end fetchUnit;

architecture SYN_Behavioral of fetchUnit is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  O : 
            out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component Mux2X1_1
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  o :
            out std_logic_vector (31 downto 0));
   end component;
   
   component InstructionRegister
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component regWithLoad32bit
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, pcToDecode_31_port, pcToDecode_30_port, 
      pcToDecode_29_port, pcToDecode_28_port, pcToDecode_27_port, 
      pcToDecode_26_port, pcToDecode_25_port, pcToDecode_24_port, 
      pcToDecode_23_port, pcToDecode_22_port, pcToDecode_21_port, 
      pcToDecode_20_port, pcToDecode_19_port, pcToDecode_18_port, 
      pcToDecode_17_port, pcToDecode_16_port, pcToDecode_15_port, 
      pcToDecode_14_port, pcToDecode_13_port, pcToDecode_12_port, 
      pcToDecode_11_port, pcToDecode_10_port, pcToDecode_9_port, 
      pcToDecode_8_port, pcToDecode_7_port, pcToDecode_6_port, 
      pcToDecode_5_port, pcToDecode_4_port, pcToDecode_3_port, 
      pcToDecode_2_port, pcToDecode_1_port, pcToDecode_0_port, 
      fromMuxToPc_31_port, fromMuxToPc_30_port, fromMuxToPc_29_port, 
      fromMuxToPc_28_port, fromMuxToPc_27_port, fromMuxToPc_26_port, 
      fromMuxToPc_25_port, fromMuxToPc_24_port, fromMuxToPc_23_port, 
      fromMuxToPc_22_port, fromMuxToPc_21_port, fromMuxToPc_20_port, 
      fromMuxToPc_19_port, fromMuxToPc_18_port, fromMuxToPc_17_port, 
      fromMuxToPc_16_port, fromMuxToPc_15_port, fromMuxToPc_14_port, 
      fromMuxToPc_13_port, fromMuxToPc_12_port, fromMuxToPc_11_port, 
      fromMuxToPc_10_port, fromMuxToPc_9_port, fromMuxToPc_8_port, 
      fromMuxToPc_7_port, fromMuxToPc_6_port, fromMuxToPc_5_port, 
      fromMuxToPc_4_port, fromMuxToPc_3_port, fromMuxToPc_2_port, 
      fromMuxToPc_1_port, fromMuxToPc_0_port, fromAdderToMux_31_port, 
      fromAdderToMux_30_port, fromAdderToMux_29_port, fromAdderToMux_28_port, 
      fromAdderToMux_27_port, fromAdderToMux_26_port, fromAdderToMux_25_port, 
      fromAdderToMux_24_port, fromAdderToMux_23_port, fromAdderToMux_22_port, 
      fromAdderToMux_21_port, fromAdderToMux_20_port, fromAdderToMux_19_port, 
      fromAdderToMux_18_port, fromAdderToMux_17_port, fromAdderToMux_16_port, 
      fromAdderToMux_15_port, fromAdderToMux_14_port, fromAdderToMux_13_port, 
      fromAdderToMux_12_port, fromAdderToMux_11_port, fromAdderToMux_10_port, 
      fromAdderToMux_9_port, fromAdderToMux_8_port, fromAdderToMux_7_port, 
      fromAdderToMux_6_port, fromAdderToMux_5_port, fromAdderToMux_4_port, 
      fromAdderToMux_3_port, fromAdderToMux_2_port, fromAdderToMux_1_port, 
      fromAdderToMux_0_port, net2804, n3 : std_logic;

begin
   PcToInstructionMemory <= ( pcToDecode_31_port, pcToDecode_30_port, 
      pcToDecode_29_port, pcToDecode_28_port, pcToDecode_27_port, 
      pcToDecode_26_port, pcToDecode_25_port, pcToDecode_24_port, 
      pcToDecode_23_port, pcToDecode_22_port, pcToDecode_21_port, 
      pcToDecode_20_port, pcToDecode_19_port, pcToDecode_18_port, 
      pcToDecode_17_port, pcToDecode_16_port, pcToDecode_15_port, 
      pcToDecode_14_port, pcToDecode_13_port, pcToDecode_12_port, 
      pcToDecode_11_port, pcToDecode_10_port, pcToDecode_9_port, 
      pcToDecode_8_port, pcToDecode_7_port, pcToDecode_6_port, 
      pcToDecode_5_port, pcToDecode_4_port, pcToDecode_3_port, 
      pcToDecode_2_port, pcToDecode_1_port, pcToDecode_0_port );
   pcToDecode <= ( pcToDecode_31_port, pcToDecode_30_port, pcToDecode_29_port, 
      pcToDecode_28_port, pcToDecode_27_port, pcToDecode_26_port, 
      pcToDecode_25_port, pcToDecode_24_port, pcToDecode_23_port, 
      pcToDecode_22_port, pcToDecode_21_port, pcToDecode_20_port, 
      pcToDecode_19_port, pcToDecode_18_port, pcToDecode_17_port, 
      pcToDecode_16_port, pcToDecode_15_port, pcToDecode_14_port, 
      pcToDecode_13_port, pcToDecode_12_port, pcToDecode_11_port, 
      pcToDecode_10_port, pcToDecode_9_port, pcToDecode_8_port, 
      pcToDecode_7_port, pcToDecode_6_port, pcToDecode_5_port, 
      pcToDecode_4_port, pcToDecode_3_port, pcToDecode_2_port, 
      pcToDecode_1_port, pcToDecode_0_port );
   
   X_Logic0_port <= '0';
   PC : regWithLoad32bit port map( clock => n3, reset => reset, load => en0, 
                           i(31) => fromMuxToPc_31_port, i(30) => 
                           fromMuxToPc_30_port, i(29) => fromMuxToPc_29_port, 
                           i(28) => fromMuxToPc_28_port, i(27) => 
                           fromMuxToPc_27_port, i(26) => fromMuxToPc_26_port, 
                           i(25) => fromMuxToPc_25_port, i(24) => 
                           fromMuxToPc_24_port, i(23) => fromMuxToPc_23_port, 
                           i(22) => fromMuxToPc_22_port, i(21) => 
                           fromMuxToPc_21_port, i(20) => fromMuxToPc_20_port, 
                           i(19) => fromMuxToPc_19_port, i(18) => 
                           fromMuxToPc_18_port, i(17) => fromMuxToPc_17_port, 
                           i(16) => fromMuxToPc_16_port, i(15) => 
                           fromMuxToPc_15_port, i(14) => fromMuxToPc_14_port, 
                           i(13) => fromMuxToPc_13_port, i(12) => 
                           fromMuxToPc_12_port, i(11) => fromMuxToPc_11_port, 
                           i(10) => fromMuxToPc_10_port, i(9) => 
                           fromMuxToPc_9_port, i(8) => fromMuxToPc_8_port, i(7)
                           => fromMuxToPc_7_port, i(6) => fromMuxToPc_6_port, 
                           i(5) => fromMuxToPc_5_port, i(4) => 
                           fromMuxToPc_4_port, i(3) => fromMuxToPc_3_port, i(2)
                           => fromMuxToPc_2_port, i(1) => fromMuxToPc_1_port, 
                           i(0) => fromMuxToPc_0_port, o(31) => 
                           pcToDecode_31_port, o(30) => pcToDecode_30_port, 
                           o(29) => pcToDecode_29_port, o(28) => 
                           pcToDecode_28_port, o(27) => pcToDecode_27_port, 
                           o(26) => pcToDecode_26_port, o(25) => 
                           pcToDecode_25_port, o(24) => pcToDecode_24_port, 
                           o(23) => pcToDecode_23_port, o(22) => 
                           pcToDecode_22_port, o(21) => pcToDecode_21_port, 
                           o(20) => pcToDecode_20_port, o(19) => 
                           pcToDecode_19_port, o(18) => pcToDecode_18_port, 
                           o(17) => pcToDecode_17_port, o(16) => 
                           pcToDecode_16_port, o(15) => pcToDecode_15_port, 
                           o(14) => pcToDecode_14_port, o(13) => 
                           pcToDecode_13_port, o(12) => pcToDecode_12_port, 
                           o(11) => pcToDecode_11_port, o(10) => 
                           pcToDecode_10_port, o(9) => pcToDecode_9_port, o(8) 
                           => pcToDecode_8_port, o(7) => pcToDecode_7_port, 
                           o(6) => pcToDecode_6_port, o(5) => pcToDecode_5_port
                           , o(4) => pcToDecode_4_port, o(3) => 
                           pcToDecode_3_port, o(2) => pcToDecode_2_port, o(1) 
                           => pcToDecode_1_port, o(0) => pcToDecode_0_port);
   IR : InstructionRegister port map( clock => n3, reset => reset, load => en0,
                           i(31) => fromInstructionMemory(31), i(30) => 
                           fromInstructionMemory(30), i(29) => 
                           fromInstructionMemory(29), i(28) => 
                           fromInstructionMemory(28), i(27) => 
                           fromInstructionMemory(27), i(26) => 
                           fromInstructionMemory(26), i(25) => 
                           fromInstructionMemory(25), i(24) => 
                           fromInstructionMemory(24), i(23) => 
                           fromInstructionMemory(23), i(22) => 
                           fromInstructionMemory(22), i(21) => 
                           fromInstructionMemory(21), i(20) => 
                           fromInstructionMemory(20), i(19) => 
                           fromInstructionMemory(19), i(18) => 
                           fromInstructionMemory(18), i(17) => 
                           fromInstructionMemory(17), i(16) => 
                           fromInstructionMemory(16), i(15) => 
                           fromInstructionMemory(15), i(14) => 
                           fromInstructionMemory(14), i(13) => 
                           fromInstructionMemory(13), i(12) => 
                           fromInstructionMemory(12), i(11) => 
                           fromInstructionMemory(11), i(10) => 
                           fromInstructionMemory(10), i(9) => 
                           fromInstructionMemory(9), i(8) => 
                           fromInstructionMemory(8), i(7) => 
                           fromInstructionMemory(7), i(6) => 
                           fromInstructionMemory(6), i(5) => 
                           fromInstructionMemory(5), i(4) => 
                           fromInstructionMemory(4), i(3) => 
                           fromInstructionMemory(3), i(2) => 
                           fromInstructionMemory(2), i(1) => 
                           fromInstructionMemory(1), i(0) => 
                           fromInstructionMemory(0), o(31) => 
                           InstructionToDecode(31), o(30) => 
                           InstructionToDecode(30), o(29) => 
                           InstructionToDecode(29), o(28) => 
                           InstructionToDecode(28), o(27) => 
                           InstructionToDecode(27), o(26) => 
                           InstructionToDecode(26), o(25) => 
                           InstructionToDecode(25), o(24) => 
                           InstructionToDecode(24), o(23) => 
                           InstructionToDecode(23), o(22) => 
                           InstructionToDecode(22), o(21) => 
                           InstructionToDecode(21), o(20) => 
                           InstructionToDecode(20), o(19) => 
                           InstructionToDecode(19), o(18) => 
                           InstructionToDecode(18), o(17) => 
                           InstructionToDecode(17), o(16) => 
                           InstructionToDecode(16), o(15) => 
                           InstructionToDecode(15), o(14) => 
                           InstructionToDecode(14), o(13) => 
                           InstructionToDecode(13), o(12) => 
                           InstructionToDecode(12), o(11) => 
                           InstructionToDecode(11), o(10) => 
                           InstructionToDecode(10), o(9) => 
                           InstructionToDecode(9), o(8) => 
                           InstructionToDecode(8), o(7) => 
                           InstructionToDecode(7), o(6) => 
                           InstructionToDecode(6), o(5) => 
                           InstructionToDecode(5), o(4) => 
                           InstructionToDecode(4), o(3) => 
                           InstructionToDecode(3), o(2) => 
                           InstructionToDecode(2), o(1) => 
                           InstructionToDecode(1), o(0) => 
                           InstructionToDecode(0));
   MUX : Mux2X1_1 port map( a(31) => next_PC(31), a(30) => next_PC(30), a(29) 
                           => next_PC(29), a(28) => next_PC(28), a(27) => 
                           next_PC(27), a(26) => next_PC(26), a(25) => 
                           next_PC(25), a(24) => next_PC(24), a(23) => 
                           next_PC(23), a(22) => next_PC(22), a(21) => 
                           next_PC(21), a(20) => next_PC(20), a(19) => 
                           next_PC(19), a(18) => next_PC(18), a(17) => 
                           next_PC(17), a(16) => next_PC(16), a(15) => 
                           next_PC(15), a(14) => next_PC(14), a(13) => 
                           next_PC(13), a(12) => next_PC(12), a(11) => 
                           next_PC(11), a(10) => next_PC(10), a(9) => 
                           next_PC(9), a(8) => next_PC(8), a(7) => next_PC(7), 
                           a(6) => next_PC(6), a(5) => next_PC(5), a(4) => 
                           next_PC(4), a(3) => next_PC(3), a(2) => next_PC(2), 
                           a(1) => next_PC(1), a(0) => next_PC(0), b(31) => 
                           fromAdderToMux_31_port, b(30) => 
                           fromAdderToMux_30_port, b(29) => 
                           fromAdderToMux_29_port, b(28) => 
                           fromAdderToMux_28_port, b(27) => 
                           fromAdderToMux_27_port, b(26) => 
                           fromAdderToMux_26_port, b(25) => 
                           fromAdderToMux_25_port, b(24) => 
                           fromAdderToMux_24_port, b(23) => 
                           fromAdderToMux_23_port, b(22) => 
                           fromAdderToMux_22_port, b(21) => 
                           fromAdderToMux_21_port, b(20) => 
                           fromAdderToMux_20_port, b(19) => 
                           fromAdderToMux_19_port, b(18) => 
                           fromAdderToMux_18_port, b(17) => 
                           fromAdderToMux_17_port, b(16) => 
                           fromAdderToMux_16_port, b(15) => 
                           fromAdderToMux_15_port, b(14) => 
                           fromAdderToMux_14_port, b(13) => 
                           fromAdderToMux_13_port, b(12) => 
                           fromAdderToMux_12_port, b(11) => 
                           fromAdderToMux_11_port, b(10) => 
                           fromAdderToMux_10_port, b(9) => 
                           fromAdderToMux_9_port, b(8) => fromAdderToMux_8_port
                           , b(7) => fromAdderToMux_7_port, b(6) => 
                           fromAdderToMux_6_port, b(5) => fromAdderToMux_5_port
                           , b(4) => fromAdderToMux_4_port, b(3) => 
                           fromAdderToMux_3_port, b(2) => fromAdderToMux_2_port
                           , b(1) => fromAdderToMux_1_port, b(0) => 
                           fromAdderToMux_0_port, sel => sel0, o(31) => 
                           fromMuxToPc_31_port, o(30) => fromMuxToPc_30_port, 
                           o(29) => fromMuxToPc_29_port, o(28) => 
                           fromMuxToPc_28_port, o(27) => fromMuxToPc_27_port, 
                           o(26) => fromMuxToPc_26_port, o(25) => 
                           fromMuxToPc_25_port, o(24) => fromMuxToPc_24_port, 
                           o(23) => fromMuxToPc_23_port, o(22) => 
                           fromMuxToPc_22_port, o(21) => fromMuxToPc_21_port, 
                           o(20) => fromMuxToPc_20_port, o(19) => 
                           fromMuxToPc_19_port, o(18) => fromMuxToPc_18_port, 
                           o(17) => fromMuxToPc_17_port, o(16) => 
                           fromMuxToPc_16_port, o(15) => fromMuxToPc_15_port, 
                           o(14) => fromMuxToPc_14_port, o(13) => 
                           fromMuxToPc_13_port, o(12) => fromMuxToPc_12_port, 
                           o(11) => fromMuxToPc_11_port, o(10) => 
                           fromMuxToPc_10_port, o(9) => fromMuxToPc_9_port, 
                           o(8) => fromMuxToPc_8_port, o(7) => 
                           fromMuxToPc_7_port, o(6) => fromMuxToPc_6_port, o(5)
                           => fromMuxToPc_5_port, o(4) => fromMuxToPc_4_port, 
                           o(3) => fromMuxToPc_3_port, o(2) => 
                           fromMuxToPc_2_port, o(1) => fromMuxToPc_1_port, o(0)
                           => fromMuxToPc_0_port);
   A : Adder port map( A(31) => pcToDecode_31_port, A(30) => pcToDecode_30_port
                           , A(29) => pcToDecode_29_port, A(28) => 
                           pcToDecode_28_port, A(27) => pcToDecode_27_port, 
                           A(26) => pcToDecode_26_port, A(25) => 
                           pcToDecode_25_port, A(24) => pcToDecode_24_port, 
                           A(23) => pcToDecode_23_port, A(22) => 
                           pcToDecode_22_port, A(21) => pcToDecode_21_port, 
                           A(20) => pcToDecode_20_port, A(19) => 
                           pcToDecode_19_port, A(18) => pcToDecode_18_port, 
                           A(17) => pcToDecode_17_port, A(16) => 
                           pcToDecode_16_port, A(15) => pcToDecode_15_port, 
                           A(14) => pcToDecode_14_port, A(13) => 
                           pcToDecode_13_port, A(12) => pcToDecode_12_port, 
                           A(11) => pcToDecode_11_port, A(10) => 
                           pcToDecode_10_port, A(9) => pcToDecode_9_port, A(8) 
                           => pcToDecode_8_port, A(7) => pcToDecode_7_port, 
                           A(6) => pcToDecode_6_port, A(5) => pcToDecode_5_port
                           , A(4) => pcToDecode_4_port, A(3) => 
                           pcToDecode_3_port, A(2) => pcToDecode_2_port, A(1) 
                           => pcToDecode_1_port, A(0) => pcToDecode_0_port, 
                           B(31) => X_Logic0_port, B(30) => X_Logic0_port, 
                           B(29) => X_Logic0_port, B(28) => X_Logic0_port, 
                           B(27) => X_Logic0_port, B(26) => X_Logic0_port, 
                           B(25) => X_Logic0_port, B(24) => X_Logic0_port, 
                           B(23) => X_Logic0_port, B(22) => X_Logic0_port, 
                           B(21) => X_Logic0_port, B(20) => X_Logic0_port, 
                           B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
                           B(17) => X_Logic0_port, B(16) => X_Logic0_port, 
                           B(15) => X_Logic0_port, B(14) => X_Logic0_port, 
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, CI => 
                           X_Logic0_port, O(31) => fromAdderToMux_31_port, 
                           O(30) => fromAdderToMux_30_port, O(29) => 
                           fromAdderToMux_29_port, O(28) => 
                           fromAdderToMux_28_port, O(27) => 
                           fromAdderToMux_27_port, O(26) => 
                           fromAdderToMux_26_port, O(25) => 
                           fromAdderToMux_25_port, O(24) => 
                           fromAdderToMux_24_port, O(23) => 
                           fromAdderToMux_23_port, O(22) => 
                           fromAdderToMux_22_port, O(21) => 
                           fromAdderToMux_21_port, O(20) => 
                           fromAdderToMux_20_port, O(19) => 
                           fromAdderToMux_19_port, O(18) => 
                           fromAdderToMux_18_port, O(17) => 
                           fromAdderToMux_17_port, O(16) => 
                           fromAdderToMux_16_port, O(15) => 
                           fromAdderToMux_15_port, O(14) => 
                           fromAdderToMux_14_port, O(13) => 
                           fromAdderToMux_13_port, O(12) => 
                           fromAdderToMux_12_port, O(11) => 
                           fromAdderToMux_11_port, O(10) => 
                           fromAdderToMux_10_port, O(9) => 
                           fromAdderToMux_9_port, O(8) => fromAdderToMux_8_port
                           , O(7) => fromAdderToMux_7_port, O(6) => 
                           fromAdderToMux_6_port, O(5) => fromAdderToMux_5_port
                           , O(4) => fromAdderToMux_4_port, O(3) => 
                           fromAdderToMux_3_port, O(2) => fromAdderToMux_2_port
                           , O(1) => fromAdderToMux_1_port, O(0) => 
                           fromAdderToMux_0_port, CO => net2804);
   U2 : BUF_X1 port map( A => clock, Z => n3);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity decodeUnit is

   port( clock, reset, en1, read_enable_portA, read_enable_portB, 
         write_enable_portW : in std_logic;  instructionWord : in 
         std_logic_vector (31 downto 0);  ID_EX_MemRead : in std_logic;  
         ID_EX_RT_Address : in std_logic_vector (4 downto 0);  writeData : in 
         std_logic_vector (31 downto 0);  writeAddress : in std_logic_vector (4
         downto 0);  pc : in std_logic_vector (31 downto 0);  sel_ext, 
         multi_cycle_operation : in std_logic;  enable_signal_PC_IF_ID, 
         selectNop : out std_logic;  outRT, outRD, outRS : out std_logic_vector
         (4 downto 0);  outIMM, outPC, outA, outB : out std_logic_vector (31 
         downto 0));

end decodeUnit;

architecture SYN_Structural of decodeUnit is

   component Mux2X1_2
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  o :
            out std_logic_vector (31 downto 0));
   end component;
   
   component extensionModule26bit
      port( i : in std_logic_vector (25 downto 0);  o : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component extensionModule
      port( i : in std_logic_vector (15 downto 0);  o : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component register_file
      port( data_in_port_w : in std_logic_vector (31 downto 0);  
            data_out_port_a, data_out_port_b : out std_logic_vector (31 downto 
            0);  address_port_a, address_port_b, address_port_w : in 
            std_logic_vector (4 downto 0);  r_signal_port_a, r_signal_port_b, 
            w_signal, reset, enable : in std_logic);
   end component;
   
   component hazardUnit
      port( RS_address, RT_address, RT_address_ID_EX : in std_logic_vector (4 
            downto 0);  MemRead_ID_EX, multi_cycle_operation : in std_logic;  
            enable_signal, sel1 : out std_logic);
   end component;
   
   component regWithEnable_5bit_1
      port( input : in std_logic_vector (4 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (4 downto 0));
   end component;
   
   component regWithEnable_5bit_2
      port( input : in std_logic_vector (4 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (4 downto 0));
   end component;
   
   component regWithEnable_5bit_3
      port( input : in std_logic_vector (4 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (4 downto 0));
   end component;
   
   component regWithEnable_1
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component regWithEnable_2
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component regWithEnable_3
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component regWithEnable_4
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   signal fromPortAToRegA_31_port, fromPortAToRegA_30_port, 
      fromPortAToRegA_29_port, fromPortAToRegA_28_port, fromPortAToRegA_27_port
      , fromPortAToRegA_26_port, fromPortAToRegA_25_port, 
      fromPortAToRegA_24_port, fromPortAToRegA_23_port, fromPortAToRegA_22_port
      , fromPortAToRegA_21_port, fromPortAToRegA_20_port, 
      fromPortAToRegA_19_port, fromPortAToRegA_18_port, fromPortAToRegA_17_port
      , fromPortAToRegA_16_port, fromPortAToRegA_15_port, 
      fromPortAToRegA_14_port, fromPortAToRegA_13_port, fromPortAToRegA_12_port
      , fromPortAToRegA_11_port, fromPortAToRegA_10_port, 
      fromPortAToRegA_9_port, fromPortAToRegA_8_port, fromPortAToRegA_7_port, 
      fromPortAToRegA_6_port, fromPortAToRegA_5_port, fromPortAToRegA_4_port, 
      fromPortAToRegA_3_port, fromPortAToRegA_2_port, fromPortAToRegA_1_port, 
      fromPortAToRegA_0_port, fromPortBToRegB_31_port, fromPortBToRegB_30_port,
      fromPortBToRegB_29_port, fromPortBToRegB_28_port, fromPortBToRegB_27_port
      , fromPortBToRegB_26_port, fromPortBToRegB_25_port, 
      fromPortBToRegB_24_port, fromPortBToRegB_23_port, fromPortBToRegB_22_port
      , fromPortBToRegB_21_port, fromPortBToRegB_20_port, 
      fromPortBToRegB_19_port, fromPortBToRegB_18_port, fromPortBToRegB_17_port
      , fromPortBToRegB_16_port, fromPortBToRegB_15_port, 
      fromPortBToRegB_14_port, fromPortBToRegB_13_port, fromPortBToRegB_12_port
      , fromPortBToRegB_11_port, fromPortBToRegB_10_port, 
      fromPortBToRegB_9_port, fromPortBToRegB_8_port, fromPortBToRegB_7_port, 
      fromPortBToRegB_6_port, fromPortBToRegB_5_port, fromPortBToRegB_4_port, 
      fromPortBToRegB_3_port, fromPortBToRegB_2_port, fromPortBToRegB_1_port, 
      fromPortBToRegB_0_port, fromFirstExtToImm_31_port, 
      fromFirstExtToImm_30_port, fromFirstExtToImm_29_port, 
      fromFirstExtToImm_28_port, fromFirstExtToImm_27_port, 
      fromFirstExtToImm_26_port, fromFirstExtToImm_25_port, 
      fromFirstExtToImm_24_port, fromFirstExtToImm_23_port, 
      fromFirstExtToImm_22_port, fromFirstExtToImm_21_port, 
      fromFirstExtToImm_20_port, fromFirstExtToImm_19_port, 
      fromFirstExtToImm_18_port, fromFirstExtToImm_17_port, 
      fromFirstExtToImm_16_port, fromFirstExtToImm_15_port, 
      fromFirstExtToImm_14_port, fromFirstExtToImm_13_port, 
      fromFirstExtToImm_12_port, fromFirstExtToImm_11_port, 
      fromFirstExtToImm_10_port, fromFirstExtToImm_9_port, 
      fromFirstExtToImm_8_port, fromFirstExtToImm_7_port, 
      fromFirstExtToImm_6_port, fromFirstExtToImm_5_port, 
      fromFirstExtToImm_4_port, fromFirstExtToImm_3_port, 
      fromFirstExtToImm_2_port, fromFirstExtToImm_1_port, 
      fromFirstExtToImm_0_port, fromSecExtToImm_31_port, 
      fromSecExtToImm_30_port, fromSecExtToImm_29_port, fromSecExtToImm_28_port
      , fromSecExtToImm_27_port, fromSecExtToImm_26_port, 
      fromSecExtToImm_25_port, fromSecExtToImm_24_port, fromSecExtToImm_23_port
      , fromSecExtToImm_22_port, fromSecExtToImm_21_port, 
      fromSecExtToImm_20_port, fromSecExtToImm_19_port, fromSecExtToImm_18_port
      , fromSecExtToImm_17_port, fromSecExtToImm_16_port, 
      fromSecExtToImm_15_port, fromSecExtToImm_14_port, fromSecExtToImm_13_port
      , fromSecExtToImm_12_port, fromSecExtToImm_11_port, 
      fromSecExtToImm_10_port, fromSecExtToImm_9_port, fromSecExtToImm_8_port, 
      fromSecExtToImm_7_port, fromSecExtToImm_6_port, fromSecExtToImm_5_port, 
      fromSecExtToImm_4_port, fromSecExtToImm_3_port, fromSecExtToImm_2_port, 
      fromSecExtToImm_1_port, fromSecExtToImm_0_port, fromMuxToImm_9_port, 
      fromMuxToImm_8_port, fromMuxToImm_7_port, fromMuxToImm_6_port, 
      fromMuxToImm_5_port, fromMuxToImm_4_port, fromMuxToImm_3_port, 
      fromMuxToImm_31_port, fromMuxToImm_30_port, fromMuxToImm_2_port, 
      fromMuxToImm_29_port, fromMuxToImm_28_port, fromMuxToImm_27_port, 
      fromMuxToImm_26_port, fromMuxToImm_25_port, fromMuxToImm_24_port, 
      fromMuxToImm_23_port, fromMuxToImm_22_port, fromMuxToImm_21_port, 
      fromMuxToImm_20_port, fromMuxToImm_1_port, fromMuxToImm_19_port, 
      fromMuxToImm_18_port, fromMuxToImm_17_port, fromMuxToImm_16_port, 
      fromMuxToImm_15_port, fromMuxToImm_14_port, fromMuxToImm_13_port, 
      fromMuxToImm_12_port, fromMuxToImm_11_port, fromMuxToImm_10_port, 
      fromMuxToImm_0_port : std_logic;

begin
   
   IMM : regWithEnable_4 port map( input(31) => fromMuxToImm_31_port, input(30)
                           => fromMuxToImm_30_port, input(29) => 
                           fromMuxToImm_29_port, input(28) => 
                           fromMuxToImm_28_port, input(27) => 
                           fromMuxToImm_27_port, input(26) => 
                           fromMuxToImm_26_port, input(25) => 
                           fromMuxToImm_25_port, input(24) => 
                           fromMuxToImm_24_port, input(23) => 
                           fromMuxToImm_23_port, input(22) => 
                           fromMuxToImm_22_port, input(21) => 
                           fromMuxToImm_21_port, input(20) => 
                           fromMuxToImm_20_port, input(19) => 
                           fromMuxToImm_19_port, input(18) => 
                           fromMuxToImm_18_port, input(17) => 
                           fromMuxToImm_17_port, input(16) => 
                           fromMuxToImm_16_port, input(15) => 
                           fromMuxToImm_15_port, input(14) => 
                           fromMuxToImm_14_port, input(13) => 
                           fromMuxToImm_13_port, input(12) => 
                           fromMuxToImm_12_port, input(11) => 
                           fromMuxToImm_11_port, input(10) => 
                           fromMuxToImm_10_port, input(9) => 
                           fromMuxToImm_9_port, input(8) => fromMuxToImm_8_port
                           , input(7) => fromMuxToImm_7_port, input(6) => 
                           fromMuxToImm_6_port, input(5) => fromMuxToImm_5_port
                           , input(4) => fromMuxToImm_4_port, input(3) => 
                           fromMuxToImm_3_port, input(2) => fromMuxToImm_2_port
                           , input(1) => fromMuxToImm_1_port, input(0) => 
                           fromMuxToImm_0_port, en => en1, clock => clock, 
                           reset => reset, output(31) => outIMM(31), output(30)
                           => outIMM(30), output(29) => outIMM(29), output(28) 
                           => outIMM(28), output(27) => outIMM(27), output(26) 
                           => outIMM(26), output(25) => outIMM(25), output(24) 
                           => outIMM(24), output(23) => outIMM(23), output(22) 
                           => outIMM(22), output(21) => outIMM(21), output(20) 
                           => outIMM(20), output(19) => outIMM(19), output(18) 
                           => outIMM(18), output(17) => outIMM(17), output(16) 
                           => outIMM(16), output(15) => outIMM(15), output(14) 
                           => outIMM(14), output(13) => outIMM(13), output(12) 
                           => outIMM(12), output(11) => outIMM(11), output(10) 
                           => outIMM(10), output(9) => outIMM(9), output(8) => 
                           outIMM(8), output(7) => outIMM(7), output(6) => 
                           outIMM(6), output(5) => outIMM(5), output(4) => 
                           outIMM(4), output(3) => outIMM(3), output(2) => 
                           outIMM(2), output(1) => outIMM(1), output(0) => 
                           outIMM(0));
   PC_R : regWithEnable_3 port map( input(31) => pc(31), input(30) => pc(30), 
                           input(29) => pc(29), input(28) => pc(28), input(27) 
                           => pc(27), input(26) => pc(26), input(25) => pc(25),
                           input(24) => pc(24), input(23) => pc(23), input(22) 
                           => pc(22), input(21) => pc(21), input(20) => pc(20),
                           input(19) => pc(19), input(18) => pc(18), input(17) 
                           => pc(17), input(16) => pc(16), input(15) => pc(15),
                           input(14) => pc(14), input(13) => pc(13), input(12) 
                           => pc(12), input(11) => pc(11), input(10) => pc(10),
                           input(9) => pc(9), input(8) => pc(8), input(7) => 
                           pc(7), input(6) => pc(6), input(5) => pc(5), 
                           input(4) => pc(4), input(3) => pc(3), input(2) => 
                           pc(2), input(1) => pc(1), input(0) => pc(0), en => 
                           en1, clock => clock, reset => reset, output(31) => 
                           outPC(31), output(30) => outPC(30), output(29) => 
                           outPC(29), output(28) => outPC(28), output(27) => 
                           outPC(27), output(26) => outPC(26), output(25) => 
                           outPC(25), output(24) => outPC(24), output(23) => 
                           outPC(23), output(22) => outPC(22), output(21) => 
                           outPC(21), output(20) => outPC(20), output(19) => 
                           outPC(19), output(18) => outPC(18), output(17) => 
                           outPC(17), output(16) => outPC(16), output(15) => 
                           outPC(15), output(14) => outPC(14), output(13) => 
                           outPC(13), output(12) => outPC(12), output(11) => 
                           outPC(11), output(10) => outPC(10), output(9) => 
                           outPC(9), output(8) => outPC(8), output(7) => 
                           outPC(7), output(6) => outPC(6), output(5) => 
                           outPC(5), output(4) => outPC(4), output(3) => 
                           outPC(3), output(2) => outPC(2), output(1) => 
                           outPC(1), output(0) => outPC(0));
   OP_A : regWithEnable_2 port map( input(31) => fromPortAToRegA_31_port, 
                           input(30) => fromPortAToRegA_30_port, input(29) => 
                           fromPortAToRegA_29_port, input(28) => 
                           fromPortAToRegA_28_port, input(27) => 
                           fromPortAToRegA_27_port, input(26) => 
                           fromPortAToRegA_26_port, input(25) => 
                           fromPortAToRegA_25_port, input(24) => 
                           fromPortAToRegA_24_port, input(23) => 
                           fromPortAToRegA_23_port, input(22) => 
                           fromPortAToRegA_22_port, input(21) => 
                           fromPortAToRegA_21_port, input(20) => 
                           fromPortAToRegA_20_port, input(19) => 
                           fromPortAToRegA_19_port, input(18) => 
                           fromPortAToRegA_18_port, input(17) => 
                           fromPortAToRegA_17_port, input(16) => 
                           fromPortAToRegA_16_port, input(15) => 
                           fromPortAToRegA_15_port, input(14) => 
                           fromPortAToRegA_14_port, input(13) => 
                           fromPortAToRegA_13_port, input(12) => 
                           fromPortAToRegA_12_port, input(11) => 
                           fromPortAToRegA_11_port, input(10) => 
                           fromPortAToRegA_10_port, input(9) => 
                           fromPortAToRegA_9_port, input(8) => 
                           fromPortAToRegA_8_port, input(7) => 
                           fromPortAToRegA_7_port, input(6) => 
                           fromPortAToRegA_6_port, input(5) => 
                           fromPortAToRegA_5_port, input(4) => 
                           fromPortAToRegA_4_port, input(3) => 
                           fromPortAToRegA_3_port, input(2) => 
                           fromPortAToRegA_2_port, input(1) => 
                           fromPortAToRegA_1_port, input(0) => 
                           fromPortAToRegA_0_port, en => en1, clock => clock, 
                           reset => reset, output(31) => outA(31), output(30) 
                           => outA(30), output(29) => outA(29), output(28) => 
                           outA(28), output(27) => outA(27), output(26) => 
                           outA(26), output(25) => outA(25), output(24) => 
                           outA(24), output(23) => outA(23), output(22) => 
                           outA(22), output(21) => outA(21), output(20) => 
                           outA(20), output(19) => outA(19), output(18) => 
                           outA(18), output(17) => outA(17), output(16) => 
                           outA(16), output(15) => outA(15), output(14) => 
                           outA(14), output(13) => outA(13), output(12) => 
                           outA(12), output(11) => outA(11), output(10) => 
                           outA(10), output(9) => outA(9), output(8) => outA(8)
                           , output(7) => outA(7), output(6) => outA(6), 
                           output(5) => outA(5), output(4) => outA(4), 
                           output(3) => outA(3), output(2) => outA(2), 
                           output(1) => outA(1), output(0) => outA(0));
   OP_B : regWithEnable_1 port map( input(31) => fromPortBToRegB_31_port, 
                           input(30) => fromPortBToRegB_30_port, input(29) => 
                           fromPortBToRegB_29_port, input(28) => 
                           fromPortBToRegB_28_port, input(27) => 
                           fromPortBToRegB_27_port, input(26) => 
                           fromPortBToRegB_26_port, input(25) => 
                           fromPortBToRegB_25_port, input(24) => 
                           fromPortBToRegB_24_port, input(23) => 
                           fromPortBToRegB_23_port, input(22) => 
                           fromPortBToRegB_22_port, input(21) => 
                           fromPortBToRegB_21_port, input(20) => 
                           fromPortBToRegB_20_port, input(19) => 
                           fromPortBToRegB_19_port, input(18) => 
                           fromPortBToRegB_18_port, input(17) => 
                           fromPortBToRegB_17_port, input(16) => 
                           fromPortBToRegB_16_port, input(15) => 
                           fromPortBToRegB_15_port, input(14) => 
                           fromPortBToRegB_14_port, input(13) => 
                           fromPortBToRegB_13_port, input(12) => 
                           fromPortBToRegB_12_port, input(11) => 
                           fromPortBToRegB_11_port, input(10) => 
                           fromPortBToRegB_10_port, input(9) => 
                           fromPortBToRegB_9_port, input(8) => 
                           fromPortBToRegB_8_port, input(7) => 
                           fromPortBToRegB_7_port, input(6) => 
                           fromPortBToRegB_6_port, input(5) => 
                           fromPortBToRegB_5_port, input(4) => 
                           fromPortBToRegB_4_port, input(3) => 
                           fromPortBToRegB_3_port, input(2) => 
                           fromPortBToRegB_2_port, input(1) => 
                           fromPortBToRegB_1_port, input(0) => 
                           fromPortBToRegB_0_port, en => en1, clock => clock, 
                           reset => reset, output(31) => outB(31), output(30) 
                           => outB(30), output(29) => outB(29), output(28) => 
                           outB(28), output(27) => outB(27), output(26) => 
                           outB(26), output(25) => outB(25), output(24) => 
                           outB(24), output(23) => outB(23), output(22) => 
                           outB(22), output(21) => outB(21), output(20) => 
                           outB(20), output(19) => outB(19), output(18) => 
                           outB(18), output(17) => outB(17), output(16) => 
                           outB(16), output(15) => outB(15), output(14) => 
                           outB(14), output(13) => outB(13), output(12) => 
                           outB(12), output(11) => outB(11), output(10) => 
                           outB(10), output(9) => outB(9), output(8) => outB(8)
                           , output(7) => outB(7), output(6) => outB(6), 
                           output(5) => outB(5), output(4) => outB(4), 
                           output(3) => outB(3), output(2) => outB(2), 
                           output(1) => outB(1), output(0) => outB(0));
   OP_RD : regWithEnable_5bit_3 port map( input(4) => instructionWord(15), 
                           input(3) => instructionWord(14), input(2) => 
                           instructionWord(13), input(1) => instructionWord(12)
                           , input(0) => instructionWord(11), en => en1, clock 
                           => clock, reset => reset, output(4) => outRD(4), 
                           output(3) => outRD(3), output(2) => outRD(2), 
                           output(1) => outRD(1), output(0) => outRD(0));
   OP_RS : regWithEnable_5bit_2 port map( input(4) => instructionWord(25), 
                           input(3) => instructionWord(24), input(2) => 
                           instructionWord(23), input(1) => instructionWord(22)
                           , input(0) => instructionWord(21), en => en1, clock 
                           => clock, reset => reset, output(4) => outRS(4), 
                           output(3) => outRS(3), output(2) => outRS(2), 
                           output(1) => outRS(1), output(0) => outRS(0));
   OP_RT : regWithEnable_5bit_1 port map( input(4) => instructionWord(20), 
                           input(3) => instructionWord(19), input(2) => 
                           instructionWord(18), input(1) => instructionWord(17)
                           , input(0) => instructionWord(16), en => en1, clock 
                           => clock, reset => reset, output(4) => outRT(4), 
                           output(3) => outRT(3), output(2) => outRT(2), 
                           output(1) => outRT(1), output(0) => outRT(0));
   HU : hazardUnit port map( RS_address(4) => instructionWord(25), 
                           RS_address(3) => instructionWord(24), RS_address(2) 
                           => instructionWord(23), RS_address(1) => 
                           instructionWord(22), RS_address(0) => 
                           instructionWord(21), RT_address(4) => 
                           instructionWord(20), RT_address(3) => 
                           instructionWord(19), RT_address(2) => 
                           instructionWord(18), RT_address(1) => 
                           instructionWord(17), RT_address(0) => 
                           instructionWord(16), RT_address_ID_EX(4) => 
                           ID_EX_RT_Address(4), RT_address_ID_EX(3) => 
                           ID_EX_RT_Address(3), RT_address_ID_EX(2) => 
                           ID_EX_RT_Address(2), RT_address_ID_EX(1) => 
                           ID_EX_RT_Address(1), RT_address_ID_EX(0) => 
                           ID_EX_RT_Address(0), MemRead_ID_EX => ID_EX_MemRead,
                           multi_cycle_operation => multi_cycle_operation, 
                           enable_signal => enable_signal_PC_IF_ID, sel1 => 
                           selectNop);
   RF : register_file port map( data_in_port_w(31) => writeData(31), 
                           data_in_port_w(30) => writeData(30), 
                           data_in_port_w(29) => writeData(29), 
                           data_in_port_w(28) => writeData(28), 
                           data_in_port_w(27) => writeData(27), 
                           data_in_port_w(26) => writeData(26), 
                           data_in_port_w(25) => writeData(25), 
                           data_in_port_w(24) => writeData(24), 
                           data_in_port_w(23) => writeData(23), 
                           data_in_port_w(22) => writeData(22), 
                           data_in_port_w(21) => writeData(21), 
                           data_in_port_w(20) => writeData(20), 
                           data_in_port_w(19) => writeData(19), 
                           data_in_port_w(18) => writeData(18), 
                           data_in_port_w(17) => writeData(17), 
                           data_in_port_w(16) => writeData(16), 
                           data_in_port_w(15) => writeData(15), 
                           data_in_port_w(14) => writeData(14), 
                           data_in_port_w(13) => writeData(13), 
                           data_in_port_w(12) => writeData(12), 
                           data_in_port_w(11) => writeData(11), 
                           data_in_port_w(10) => writeData(10), 
                           data_in_port_w(9) => writeData(9), data_in_port_w(8)
                           => writeData(8), data_in_port_w(7) => writeData(7), 
                           data_in_port_w(6) => writeData(6), data_in_port_w(5)
                           => writeData(5), data_in_port_w(4) => writeData(4), 
                           data_in_port_w(3) => writeData(3), data_in_port_w(2)
                           => writeData(2), data_in_port_w(1) => writeData(1), 
                           data_in_port_w(0) => writeData(0), 
                           data_out_port_a(31) => fromPortAToRegA_31_port, 
                           data_out_port_a(30) => fromPortAToRegA_30_port, 
                           data_out_port_a(29) => fromPortAToRegA_29_port, 
                           data_out_port_a(28) => fromPortAToRegA_28_port, 
                           data_out_port_a(27) => fromPortAToRegA_27_port, 
                           data_out_port_a(26) => fromPortAToRegA_26_port, 
                           data_out_port_a(25) => fromPortAToRegA_25_port, 
                           data_out_port_a(24) => fromPortAToRegA_24_port, 
                           data_out_port_a(23) => fromPortAToRegA_23_port, 
                           data_out_port_a(22) => fromPortAToRegA_22_port, 
                           data_out_port_a(21) => fromPortAToRegA_21_port, 
                           data_out_port_a(20) => fromPortAToRegA_20_port, 
                           data_out_port_a(19) => fromPortAToRegA_19_port, 
                           data_out_port_a(18) => fromPortAToRegA_18_port, 
                           data_out_port_a(17) => fromPortAToRegA_17_port, 
                           data_out_port_a(16) => fromPortAToRegA_16_port, 
                           data_out_port_a(15) => fromPortAToRegA_15_port, 
                           data_out_port_a(14) => fromPortAToRegA_14_port, 
                           data_out_port_a(13) => fromPortAToRegA_13_port, 
                           data_out_port_a(12) => fromPortAToRegA_12_port, 
                           data_out_port_a(11) => fromPortAToRegA_11_port, 
                           data_out_port_a(10) => fromPortAToRegA_10_port, 
                           data_out_port_a(9) => fromPortAToRegA_9_port, 
                           data_out_port_a(8) => fromPortAToRegA_8_port, 
                           data_out_port_a(7) => fromPortAToRegA_7_port, 
                           data_out_port_a(6) => fromPortAToRegA_6_port, 
                           data_out_port_a(5) => fromPortAToRegA_5_port, 
                           data_out_port_a(4) => fromPortAToRegA_4_port, 
                           data_out_port_a(3) => fromPortAToRegA_3_port, 
                           data_out_port_a(2) => fromPortAToRegA_2_port, 
                           data_out_port_a(1) => fromPortAToRegA_1_port, 
                           data_out_port_a(0) => fromPortAToRegA_0_port, 
                           data_out_port_b(31) => fromPortBToRegB_31_port, 
                           data_out_port_b(30) => fromPortBToRegB_30_port, 
                           data_out_port_b(29) => fromPortBToRegB_29_port, 
                           data_out_port_b(28) => fromPortBToRegB_28_port, 
                           data_out_port_b(27) => fromPortBToRegB_27_port, 
                           data_out_port_b(26) => fromPortBToRegB_26_port, 
                           data_out_port_b(25) => fromPortBToRegB_25_port, 
                           data_out_port_b(24) => fromPortBToRegB_24_port, 
                           data_out_port_b(23) => fromPortBToRegB_23_port, 
                           data_out_port_b(22) => fromPortBToRegB_22_port, 
                           data_out_port_b(21) => fromPortBToRegB_21_port, 
                           data_out_port_b(20) => fromPortBToRegB_20_port, 
                           data_out_port_b(19) => fromPortBToRegB_19_port, 
                           data_out_port_b(18) => fromPortBToRegB_18_port, 
                           data_out_port_b(17) => fromPortBToRegB_17_port, 
                           data_out_port_b(16) => fromPortBToRegB_16_port, 
                           data_out_port_b(15) => fromPortBToRegB_15_port, 
                           data_out_port_b(14) => fromPortBToRegB_14_port, 
                           data_out_port_b(13) => fromPortBToRegB_13_port, 
                           data_out_port_b(12) => fromPortBToRegB_12_port, 
                           data_out_port_b(11) => fromPortBToRegB_11_port, 
                           data_out_port_b(10) => fromPortBToRegB_10_port, 
                           data_out_port_b(9) => fromPortBToRegB_9_port, 
                           data_out_port_b(8) => fromPortBToRegB_8_port, 
                           data_out_port_b(7) => fromPortBToRegB_7_port, 
                           data_out_port_b(6) => fromPortBToRegB_6_port, 
                           data_out_port_b(5) => fromPortBToRegB_5_port, 
                           data_out_port_b(4) => fromPortBToRegB_4_port, 
                           data_out_port_b(3) => fromPortBToRegB_3_port, 
                           data_out_port_b(2) => fromPortBToRegB_2_port, 
                           data_out_port_b(1) => fromPortBToRegB_1_port, 
                           data_out_port_b(0) => fromPortBToRegB_0_port, 
                           address_port_a(4) => instructionWord(25), 
                           address_port_a(3) => instructionWord(24), 
                           address_port_a(2) => instructionWord(23), 
                           address_port_a(1) => instructionWord(22), 
                           address_port_a(0) => instructionWord(21), 
                           address_port_b(4) => instructionWord(20), 
                           address_port_b(3) => instructionWord(19), 
                           address_port_b(2) => instructionWord(18), 
                           address_port_b(1) => instructionWord(17), 
                           address_port_b(0) => instructionWord(16), 
                           address_port_w(4) => writeAddress(4), 
                           address_port_w(3) => writeAddress(3), 
                           address_port_w(2) => writeAddress(2), 
                           address_port_w(1) => writeAddress(1), 
                           address_port_w(0) => writeAddress(0), 
                           r_signal_port_a => read_enable_portA, 
                           r_signal_port_b => read_enable_portB, w_signal => 
                           write_enable_portW, reset => reset, enable => en1);
   EXT1 : extensionModule port map( i(15) => instructionWord(15), i(14) => 
                           instructionWord(14), i(13) => instructionWord(13), 
                           i(12) => instructionWord(12), i(11) => 
                           instructionWord(11), i(10) => instructionWord(10), 
                           i(9) => instructionWord(9), i(8) => 
                           instructionWord(8), i(7) => instructionWord(7), i(6)
                           => instructionWord(6), i(5) => instructionWord(5), 
                           i(4) => instructionWord(4), i(3) => 
                           instructionWord(3), i(2) => instructionWord(2), i(1)
                           => instructionWord(1), i(0) => instructionWord(0), 
                           o(31) => fromFirstExtToImm_31_port, o(30) => 
                           fromFirstExtToImm_30_port, o(29) => 
                           fromFirstExtToImm_29_port, o(28) => 
                           fromFirstExtToImm_28_port, o(27) => 
                           fromFirstExtToImm_27_port, o(26) => 
                           fromFirstExtToImm_26_port, o(25) => 
                           fromFirstExtToImm_25_port, o(24) => 
                           fromFirstExtToImm_24_port, o(23) => 
                           fromFirstExtToImm_23_port, o(22) => 
                           fromFirstExtToImm_22_port, o(21) => 
                           fromFirstExtToImm_21_port, o(20) => 
                           fromFirstExtToImm_20_port, o(19) => 
                           fromFirstExtToImm_19_port, o(18) => 
                           fromFirstExtToImm_18_port, o(17) => 
                           fromFirstExtToImm_17_port, o(16) => 
                           fromFirstExtToImm_16_port, o(15) => 
                           fromFirstExtToImm_15_port, o(14) => 
                           fromFirstExtToImm_14_port, o(13) => 
                           fromFirstExtToImm_13_port, o(12) => 
                           fromFirstExtToImm_12_port, o(11) => 
                           fromFirstExtToImm_11_port, o(10) => 
                           fromFirstExtToImm_10_port, o(9) => 
                           fromFirstExtToImm_9_port, o(8) => 
                           fromFirstExtToImm_8_port, o(7) => 
                           fromFirstExtToImm_7_port, o(6) => 
                           fromFirstExtToImm_6_port, o(5) => 
                           fromFirstExtToImm_5_port, o(4) => 
                           fromFirstExtToImm_4_port, o(3) => 
                           fromFirstExtToImm_3_port, o(2) => 
                           fromFirstExtToImm_2_port, o(1) => 
                           fromFirstExtToImm_1_port, o(0) => 
                           fromFirstExtToImm_0_port);
   EXT2 : extensionModule26bit port map( i(25) => instructionWord(25), i(24) =>
                           instructionWord(24), i(23) => instructionWord(23), 
                           i(22) => instructionWord(22), i(21) => 
                           instructionWord(21), i(20) => instructionWord(20), 
                           i(19) => instructionWord(19), i(18) => 
                           instructionWord(18), i(17) => instructionWord(17), 
                           i(16) => instructionWord(16), i(15) => 
                           instructionWord(15), i(14) => instructionWord(14), 
                           i(13) => instructionWord(13), i(12) => 
                           instructionWord(12), i(11) => instructionWord(11), 
                           i(10) => instructionWord(10), i(9) => 
                           instructionWord(9), i(8) => instructionWord(8), i(7)
                           => instructionWord(7), i(6) => instructionWord(6), 
                           i(5) => instructionWord(5), i(4) => 
                           instructionWord(4), i(3) => instructionWord(3), i(2)
                           => instructionWord(2), i(1) => instructionWord(1), 
                           i(0) => instructionWord(0), o(31) => 
                           fromSecExtToImm_31_port, o(30) => 
                           fromSecExtToImm_30_port, o(29) => 
                           fromSecExtToImm_29_port, o(28) => 
                           fromSecExtToImm_28_port, o(27) => 
                           fromSecExtToImm_27_port, o(26) => 
                           fromSecExtToImm_26_port, o(25) => 
                           fromSecExtToImm_25_port, o(24) => 
                           fromSecExtToImm_24_port, o(23) => 
                           fromSecExtToImm_23_port, o(22) => 
                           fromSecExtToImm_22_port, o(21) => 
                           fromSecExtToImm_21_port, o(20) => 
                           fromSecExtToImm_20_port, o(19) => 
                           fromSecExtToImm_19_port, o(18) => 
                           fromSecExtToImm_18_port, o(17) => 
                           fromSecExtToImm_17_port, o(16) => 
                           fromSecExtToImm_16_port, o(15) => 
                           fromSecExtToImm_15_port, o(14) => 
                           fromSecExtToImm_14_port, o(13) => 
                           fromSecExtToImm_13_port, o(12) => 
                           fromSecExtToImm_12_port, o(11) => 
                           fromSecExtToImm_11_port, o(10) => 
                           fromSecExtToImm_10_port, o(9) => 
                           fromSecExtToImm_9_port, o(8) => 
                           fromSecExtToImm_8_port, o(7) => 
                           fromSecExtToImm_7_port, o(6) => 
                           fromSecExtToImm_6_port, o(5) => 
                           fromSecExtToImm_5_port, o(4) => 
                           fromSecExtToImm_4_port, o(3) => 
                           fromSecExtToImm_3_port, o(2) => 
                           fromSecExtToImm_2_port, o(1) => 
                           fromSecExtToImm_1_port, o(0) => 
                           fromSecExtToImm_0_port);
   MUXEXT : Mux2X1_2 port map( a(31) => fromFirstExtToImm_31_port, a(30) => 
                           fromFirstExtToImm_30_port, a(29) => 
                           fromFirstExtToImm_29_port, a(28) => 
                           fromFirstExtToImm_28_port, a(27) => 
                           fromFirstExtToImm_27_port, a(26) => 
                           fromFirstExtToImm_26_port, a(25) => 
                           fromFirstExtToImm_25_port, a(24) => 
                           fromFirstExtToImm_24_port, a(23) => 
                           fromFirstExtToImm_23_port, a(22) => 
                           fromFirstExtToImm_22_port, a(21) => 
                           fromFirstExtToImm_21_port, a(20) => 
                           fromFirstExtToImm_20_port, a(19) => 
                           fromFirstExtToImm_19_port, a(18) => 
                           fromFirstExtToImm_18_port, a(17) => 
                           fromFirstExtToImm_17_port, a(16) => 
                           fromFirstExtToImm_16_port, a(15) => 
                           fromFirstExtToImm_15_port, a(14) => 
                           fromFirstExtToImm_14_port, a(13) => 
                           fromFirstExtToImm_13_port, a(12) => 
                           fromFirstExtToImm_12_port, a(11) => 
                           fromFirstExtToImm_11_port, a(10) => 
                           fromFirstExtToImm_10_port, a(9) => 
                           fromFirstExtToImm_9_port, a(8) => 
                           fromFirstExtToImm_8_port, a(7) => 
                           fromFirstExtToImm_7_port, a(6) => 
                           fromFirstExtToImm_6_port, a(5) => 
                           fromFirstExtToImm_5_port, a(4) => 
                           fromFirstExtToImm_4_port, a(3) => 
                           fromFirstExtToImm_3_port, a(2) => 
                           fromFirstExtToImm_2_port, a(1) => 
                           fromFirstExtToImm_1_port, a(0) => 
                           fromFirstExtToImm_0_port, b(31) => 
                           fromSecExtToImm_31_port, b(30) => 
                           fromSecExtToImm_30_port, b(29) => 
                           fromSecExtToImm_29_port, b(28) => 
                           fromSecExtToImm_28_port, b(27) => 
                           fromSecExtToImm_27_port, b(26) => 
                           fromSecExtToImm_26_port, b(25) => 
                           fromSecExtToImm_25_port, b(24) => 
                           fromSecExtToImm_24_port, b(23) => 
                           fromSecExtToImm_23_port, b(22) => 
                           fromSecExtToImm_22_port, b(21) => 
                           fromSecExtToImm_21_port, b(20) => 
                           fromSecExtToImm_20_port, b(19) => 
                           fromSecExtToImm_19_port, b(18) => 
                           fromSecExtToImm_18_port, b(17) => 
                           fromSecExtToImm_17_port, b(16) => 
                           fromSecExtToImm_16_port, b(15) => 
                           fromSecExtToImm_15_port, b(14) => 
                           fromSecExtToImm_14_port, b(13) => 
                           fromSecExtToImm_13_port, b(12) => 
                           fromSecExtToImm_12_port, b(11) => 
                           fromSecExtToImm_11_port, b(10) => 
                           fromSecExtToImm_10_port, b(9) => 
                           fromSecExtToImm_9_port, b(8) => 
                           fromSecExtToImm_8_port, b(7) => 
                           fromSecExtToImm_7_port, b(6) => 
                           fromSecExtToImm_6_port, b(5) => 
                           fromSecExtToImm_5_port, b(4) => 
                           fromSecExtToImm_4_port, b(3) => 
                           fromSecExtToImm_3_port, b(2) => 
                           fromSecExtToImm_2_port, b(1) => 
                           fromSecExtToImm_1_port, b(0) => 
                           fromSecExtToImm_0_port, sel => sel_ext, o(31) => 
                           fromMuxToImm_31_port, o(30) => fromMuxToImm_30_port,
                           o(29) => fromMuxToImm_29_port, o(28) => 
                           fromMuxToImm_28_port, o(27) => fromMuxToImm_27_port,
                           o(26) => fromMuxToImm_26_port, o(25) => 
                           fromMuxToImm_25_port, o(24) => fromMuxToImm_24_port,
                           o(23) => fromMuxToImm_23_port, o(22) => 
                           fromMuxToImm_22_port, o(21) => fromMuxToImm_21_port,
                           o(20) => fromMuxToImm_20_port, o(19) => 
                           fromMuxToImm_19_port, o(18) => fromMuxToImm_18_port,
                           o(17) => fromMuxToImm_17_port, o(16) => 
                           fromMuxToImm_16_port, o(15) => fromMuxToImm_15_port,
                           o(14) => fromMuxToImm_14_port, o(13) => 
                           fromMuxToImm_13_port, o(12) => fromMuxToImm_12_port,
                           o(11) => fromMuxToImm_11_port, o(10) => 
                           fromMuxToImm_10_port, o(9) => fromMuxToImm_9_port, 
                           o(8) => fromMuxToImm_8_port, o(7) => 
                           fromMuxToImm_7_port, o(6) => fromMuxToImm_6_port, 
                           o(5) => fromMuxToImm_5_port, o(4) => 
                           fromMuxToImm_4_port, o(3) => fromMuxToImm_3_port, 
                           o(2) => fromMuxToImm_2_port, o(1) => 
                           fromMuxToImm_1_port, o(0) => fromMuxToImm_0_port);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity executionUnit is

   port( clock, reset : in std_logic;  operand_a, operand_b, operand_imm, 
         operand_pc, forward_exe, forward_mem : in std_logic_vector (31 downto 
         0);  EX_MEM_write, MEM_WB_write : in std_logic;  MEM_WB_rd, ID_EX_Rd, 
         ID_EX_Rs, ID_EX_Rt : in std_logic_vector (4 downto 0);  enable, sel_1,
         sel_2, sel_3 : in std_logic;  func : in std_logic_vector (10 downto 0)
         ;  EX_MEM_rd : inout std_logic_vector (4 downto 0);  
         out_res_operand_one, out_res_operand_two, next_pc : out 
         std_logic_vector (31 downto 0);  jump, multi_cycle_operation : out 
         std_logic);

end executionUnit;

architecture SYN_Structural of executionUnit is

   component mux3_1_1
      port( operand_one, operand_two, operand_three : in std_logic_vector (31 
            downto 0);  sel : in std_logic_vector (1 downto 0);  out_res : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component mux3_1_0
      port( operand_one, operand_two, operand_three : in std_logic_vector (31 
            downto 0);  sel : in std_logic_vector (1 downto 0);  out_res : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component Mux2X1_3
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  o :
            out std_logic_vector (31 downto 0));
   end component;
   
   component Mux2X1_4
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  o :
            out std_logic_vector (31 downto 0));
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_8
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component pentium4_adder_XBIT32_NBIT4_0
      port( A, B : in std_logic_vector (31 downto 0);  C_0 : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component comparator
      port( A, B : in std_logic_vector (31 downto 0);  Sel : in 
            std_logic_vector (2 downto 0);  O : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_100_1
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_100_0
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_011_1
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_011_0
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_010_1
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_010_0
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_001_1
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_001_0
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_000_1
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component positive_latch_on_000_0
      port( d : in std_logic_vector (31 downto 0);  enable : in 
            std_logic_vector (2 downto 0);  q : out std_logic_vector (31 downto
            0));
   end component;
   
   component logicUnitT2_data_size32
      port( operand_a, operand_b : in std_logic_vector (31 downto 0);  type_op 
            : in std_logic_vector (3 downto 0);  result : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component mux5x1
      port( a, b, c, d, e : in std_logic_vector (31 downto 0);  enable : in 
            std_logic;  sel : in std_logic_vector (2 downto 0);  out_res : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component booths_mul_N_bit16
      port( multiplier, multiplicand : in std_logic_vector (15 downto 0);  
            product : out std_logic_vector (31 downto 0));
   end component;
   
   component Shifter_NBIT32
      port( left_right, logic_Arith, shift_rot : in std_logic;  a, b : in 
            std_logic_vector (31 downto 0);  o : out std_logic_vector (31 
            downto 0));
   end component;
   
   component regWithEnable_5
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component DIVIDER_N_op32
      port( CLK, START, RESET : in std_logic;  BUSY : out std_logic;  DIVIDEND,
            DIVISOR : in std_logic_vector (31 downto 0);  QUOTIENT, RESIDUAL : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component Mux2X1_5
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  o :
            out std_logic_vector (31 downto 0));
   end component;
   
   component forwarding_unit
      port( EX_MEM_write : in std_logic;  EX_MEM_Rd, ID_EX_Rs, ID_EX_Rt : in 
            std_logic_vector (4 downto 0);  MEM_WB_write : in std_logic;  
            MEM_WB_Rd : in std_logic_vector (4 downto 0);  sel_mux_high, 
            sel_mux_low : out std_logic_vector (1 downto 0));
   end component;
   
   component mux_2_1_5bit
      port( a, b : in std_logic_vector (4 downto 0);  sel : in std_logic;  o : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component regWithEnable_5bit_4
      port( input : in std_logic_vector (4 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (4 downto 0));
   end component;
   
   component cu_exe
      port( reset : in std_logic;  func : in std_logic_vector (10 downto 0);  
            busy_div : in std_logic;  multi_cycle_operation, enable : out 
            std_logic;  sel_signal_5X1 : out std_logic_vector (2 downto 0);  
            sel_signal_2X1, start_div : out std_logic;  cmd_t2 : out 
            std_logic_vector (3 downto 0);  carry_in, left_right, logic_Arith, 
            shift_rot : out std_logic;  sel_comparator : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component regWithEnable_6
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   signal jump_port, busy, enable_mux_4_1, sel_signal_5_1_2_port, 
      sel_signal_5_1_1_port, sel_signal_5_1_0_port, sel_signal_2_1, start_div, 
      signal_cmd_t2_3_port, signal_cmd_t2_2_port, signal_cmd_t2_1_port, 
      signal_cmd_t2_0_port, carry_in, left_right, logic_Arith, shift_rot, 
      sel_comparator_2_port, sel_comparator_1_port, sel_comparator_0_port, 
      EX_MEM_rd_next_4_port, EX_MEM_rd_next_3_port, EX_MEM_rd_next_2_port, 
      EX_MEM_rd_next_1_port, EX_MEM_rd_next_0_port, sel_mux_3_1_high_1_port, 
      sel_mux_3_1_high_0_port, sel_mux_3_1_low_1_port, sel_mux_3_1_low_0_port, 
      quotient_31_port, quotient_30_port, quotient_29_port, quotient_28_port, 
      quotient_27_port, quotient_26_port, quotient_25_port, quotient_24_port, 
      quotient_23_port, quotient_22_port, quotient_21_port, quotient_20_port, 
      quotient_19_port, quotient_18_port, quotient_17_port, quotient_16_port, 
      quotient_15_port, quotient_14_port, quotient_13_port, quotient_12_port, 
      quotient_11_port, quotient_10_port, quotient_9_port, quotient_8_port, 
      quotient_7_port, quotient_6_port, quotient_5_port, quotient_4_port, 
      quotient_3_port, quotient_2_port, quotient_1_port, quotient_0_port, 
      from_mux_4_1_to_mux_2_1_31_port, from_mux_4_1_to_mux_2_1_30_port, 
      from_mux_4_1_to_mux_2_1_29_port, from_mux_4_1_to_mux_2_1_28_port, 
      from_mux_4_1_to_mux_2_1_27_port, from_mux_4_1_to_mux_2_1_26_port, 
      from_mux_4_1_to_mux_2_1_25_port, from_mux_4_1_to_mux_2_1_24_port, 
      from_mux_4_1_to_mux_2_1_23_port, from_mux_4_1_to_mux_2_1_22_port, 
      from_mux_4_1_to_mux_2_1_21_port, from_mux_4_1_to_mux_2_1_20_port, 
      from_mux_4_1_to_mux_2_1_19_port, from_mux_4_1_to_mux_2_1_18_port, 
      from_mux_4_1_to_mux_2_1_17_port, from_mux_4_1_to_mux_2_1_16_port, 
      from_mux_4_1_to_mux_2_1_15_port, from_mux_4_1_to_mux_2_1_14_port, 
      from_mux_4_1_to_mux_2_1_13_port, from_mux_4_1_to_mux_2_1_12_port, 
      from_mux_4_1_to_mux_2_1_11_port, from_mux_4_1_to_mux_2_1_10_port, 
      from_mux_4_1_to_mux_2_1_9_port, from_mux_4_1_to_mux_2_1_8_port, 
      from_mux_4_1_to_mux_2_1_7_port, from_mux_4_1_to_mux_2_1_6_port, 
      from_mux_4_1_to_mux_2_1_5_port, from_mux_4_1_to_mux_2_1_4_port, 
      from_mux_4_1_to_mux_2_1_3_port, from_mux_4_1_to_mux_2_1_2_port, 
      from_mux_4_1_to_mux_2_1_1_port, from_mux_4_1_to_mux_2_1_0_port, 
      from_mux_2_1_to_latch_high_31_port, from_mux_2_1_to_latch_high_30_port, 
      from_mux_2_1_to_latch_high_29_port, from_mux_2_1_to_latch_high_28_port, 
      from_mux_2_1_to_latch_high_27_port, from_mux_2_1_to_latch_high_26_port, 
      from_mux_2_1_to_latch_high_25_port, from_mux_2_1_to_latch_high_24_port, 
      from_mux_2_1_to_latch_high_23_port, from_mux_2_1_to_latch_high_22_port, 
      from_mux_2_1_to_latch_high_21_port, from_mux_2_1_to_latch_high_20_port, 
      from_mux_2_1_to_latch_high_19_port, from_mux_2_1_to_latch_high_18_port, 
      from_mux_2_1_to_latch_high_17_port, from_mux_2_1_to_latch_high_16_port, 
      from_mux_2_1_to_latch_high_15_port, from_mux_2_1_to_latch_high_14_port, 
      from_mux_2_1_to_latch_high_13_port, from_mux_2_1_to_latch_high_12_port, 
      from_mux_2_1_to_latch_high_11_port, from_mux_2_1_to_latch_high_10_port, 
      from_mux_2_1_to_latch_high_9_port, from_mux_2_1_to_latch_high_8_port, 
      from_mux_2_1_to_latch_high_7_port, from_mux_2_1_to_latch_high_6_port, 
      from_mux_2_1_to_latch_high_5_port, from_mux_2_1_to_latch_high_4_port, 
      from_mux_2_1_to_latch_high_3_port, from_mux_2_1_to_latch_high_2_port, 
      from_mux_2_1_to_latch_high_1_port, from_mux_2_1_to_latch_high_0_port, 
      from_mux_2_1_to_latch_low_31_port, from_mux_2_1_to_latch_low_30_port, 
      from_mux_2_1_to_latch_low_29_port, from_mux_2_1_to_latch_low_28_port, 
      from_mux_2_1_to_latch_low_27_port, from_mux_2_1_to_latch_low_26_port, 
      from_mux_2_1_to_latch_low_25_port, from_mux_2_1_to_latch_low_24_port, 
      from_mux_2_1_to_latch_low_23_port, from_mux_2_1_to_latch_low_22_port, 
      from_mux_2_1_to_latch_low_21_port, from_mux_2_1_to_latch_low_20_port, 
      from_mux_2_1_to_latch_low_19_port, from_mux_2_1_to_latch_low_18_port, 
      from_mux_2_1_to_latch_low_17_port, from_mux_2_1_to_latch_low_16_port, 
      from_mux_2_1_to_latch_low_15_port, from_mux_2_1_to_latch_low_14_port, 
      from_mux_2_1_to_latch_low_13_port, from_mux_2_1_to_latch_low_12_port, 
      from_mux_2_1_to_latch_low_11_port, from_mux_2_1_to_latch_low_10_port, 
      from_mux_2_1_to_latch_low_9_port, from_mux_2_1_to_latch_low_8_port, 
      from_mux_2_1_to_latch_low_7_port, from_mux_2_1_to_latch_low_6_port, 
      from_mux_2_1_to_latch_low_5_port, from_mux_2_1_to_latch_low_4_port, 
      from_mux_2_1_to_latch_low_3_port, from_mux_2_1_to_latch_low_2_port, 
      from_mux_2_1_to_latch_low_1_port, from_mux_2_1_to_latch_low_0_port, 
      from_latch_to_shifter_op1_31_port, from_latch_to_shifter_op1_30_port, 
      from_latch_to_shifter_op1_29_port, from_latch_to_shifter_op1_28_port, 
      from_latch_to_shifter_op1_27_port, from_latch_to_shifter_op1_26_port, 
      from_latch_to_shifter_op1_25_port, from_latch_to_shifter_op1_24_port, 
      from_latch_to_shifter_op1_23_port, from_latch_to_shifter_op1_22_port, 
      from_latch_to_shifter_op1_21_port, from_latch_to_shifter_op1_20_port, 
      from_latch_to_shifter_op1_19_port, from_latch_to_shifter_op1_18_port, 
      from_latch_to_shifter_op1_17_port, from_latch_to_shifter_op1_16_port, 
      from_latch_to_shifter_op1_15_port, from_latch_to_shifter_op1_14_port, 
      from_latch_to_shifter_op1_13_port, from_latch_to_shifter_op1_12_port, 
      from_latch_to_shifter_op1_11_port, from_latch_to_shifter_op1_10_port, 
      from_latch_to_shifter_op1_9_port, from_latch_to_shifter_op1_8_port, 
      from_latch_to_shifter_op1_7_port, from_latch_to_shifter_op1_6_port, 
      from_latch_to_shifter_op1_5_port, from_latch_to_shifter_op1_4_port, 
      from_latch_to_shifter_op1_3_port, from_latch_to_shifter_op1_2_port, 
      from_latch_to_shifter_op1_1_port, from_latch_to_shifter_op1_0_port, 
      from_latch_to_shifter_op2_31_port, from_latch_to_shifter_op2_30_port, 
      from_latch_to_shifter_op2_29_port, from_latch_to_shifter_op2_28_port, 
      from_latch_to_shifter_op2_27_port, from_latch_to_shifter_op2_26_port, 
      from_latch_to_shifter_op2_25_port, from_latch_to_shifter_op2_24_port, 
      from_latch_to_shifter_op2_23_port, from_latch_to_shifter_op2_22_port, 
      from_latch_to_shifter_op2_21_port, from_latch_to_shifter_op2_20_port, 
      from_latch_to_shifter_op2_19_port, from_latch_to_shifter_op2_18_port, 
      from_latch_to_shifter_op2_17_port, from_latch_to_shifter_op2_16_port, 
      from_latch_to_shifter_op2_15_port, from_latch_to_shifter_op2_14_port, 
      from_latch_to_shifter_op2_13_port, from_latch_to_shifter_op2_12_port, 
      from_latch_to_shifter_op2_11_port, from_latch_to_shifter_op2_10_port, 
      from_latch_to_shifter_op2_9_port, from_latch_to_shifter_op2_8_port, 
      from_latch_to_shifter_op2_7_port, from_latch_to_shifter_op2_6_port, 
      from_latch_to_shifter_op2_5_port, from_latch_to_shifter_op2_4_port, 
      from_latch_to_shifter_op2_3_port, from_latch_to_shifter_op2_2_port, 
      from_latch_to_shifter_op2_1_port, from_latch_to_shifter_op2_0_port, 
      from_shifter_to_mux_31_port, from_shifter_to_mux_30_port, 
      from_shifter_to_mux_29_port, from_shifter_to_mux_28_port, 
      from_shifter_to_mux_27_port, from_shifter_to_mux_26_port, 
      from_shifter_to_mux_25_port, from_shifter_to_mux_24_port, 
      from_shifter_to_mux_23_port, from_shifter_to_mux_22_port, 
      from_shifter_to_mux_21_port, from_shifter_to_mux_20_port, 
      from_shifter_to_mux_19_port, from_shifter_to_mux_18_port, 
      from_shifter_to_mux_17_port, from_shifter_to_mux_16_port, 
      from_shifter_to_mux_15_port, from_shifter_to_mux_14_port, 
      from_shifter_to_mux_13_port, from_shifter_to_mux_12_port, 
      from_shifter_to_mux_11_port, from_shifter_to_mux_10_port, 
      from_shifter_to_mux_9_port, from_shifter_to_mux_8_port, 
      from_shifter_to_mux_7_port, from_shifter_to_mux_6_port, 
      from_shifter_to_mux_5_port, from_shifter_to_mux_4_port, 
      from_shifter_to_mux_3_port, from_shifter_to_mux_2_port, 
      from_shifter_to_mux_1_port, from_shifter_to_mux_0_port, 
      from_latch_to_mul_op2_15_port, from_latch_to_mul_op2_14_port, 
      from_latch_to_mul_op2_13_port, from_latch_to_mul_op2_12_port, 
      from_latch_to_mul_op2_11_port, from_latch_to_mul_op2_10_port, 
      from_latch_to_mul_op2_9_port, from_latch_to_mul_op2_8_port, 
      from_latch_to_mul_op2_7_port, from_latch_to_mul_op2_6_port, 
      from_latch_to_mul_op2_5_port, from_latch_to_mul_op2_4_port, 
      from_latch_to_mul_op2_3_port, from_latch_to_mul_op2_2_port, 
      from_latch_to_mul_op2_1_port, from_latch_to_mul_op2_0_port, 
      from_latch_to_mul_op1_15_port, from_latch_to_mul_op1_14_port, 
      from_latch_to_mul_op1_13_port, from_latch_to_mul_op1_12_port, 
      from_latch_to_mul_op1_11_port, from_latch_to_mul_op1_10_port, 
      from_latch_to_mul_op1_9_port, from_latch_to_mul_op1_8_port, 
      from_latch_to_mul_op1_7_port, from_latch_to_mul_op1_6_port, 
      from_latch_to_mul_op1_5_port, from_latch_to_mul_op1_4_port, 
      from_latch_to_mul_op1_3_port, from_latch_to_mul_op1_2_port, 
      from_latch_to_mul_op1_1_port, from_latch_to_mul_op1_0_port, 
      from_mul_to_mux_31_port, from_mul_to_mux_30_port, from_mul_to_mux_29_port
      , from_mul_to_mux_28_port, from_mul_to_mux_27_port, 
      from_mul_to_mux_26_port, from_mul_to_mux_25_port, from_mul_to_mux_24_port
      , from_mul_to_mux_23_port, from_mul_to_mux_22_port, 
      from_mul_to_mux_21_port, from_mul_to_mux_20_port, from_mul_to_mux_19_port
      , from_mul_to_mux_18_port, from_mul_to_mux_17_port, 
      from_mul_to_mux_16_port, from_mul_to_mux_15_port, from_mul_to_mux_14_port
      , from_mul_to_mux_13_port, from_mul_to_mux_12_port, 
      from_mul_to_mux_11_port, from_mul_to_mux_10_port, from_mul_to_mux_9_port,
      from_mul_to_mux_8_port, from_mul_to_mux_7_port, from_mul_to_mux_6_port, 
      from_mul_to_mux_5_port, from_mul_to_mux_4_port, from_mul_to_mux_3_port, 
      from_mul_to_mux_2_port, from_mul_to_mux_1_port, from_mul_to_mux_0_port, 
      from_adder_to_mux_31_port, from_adder_to_mux_30_port, 
      from_adder_to_mux_29_port, from_adder_to_mux_28_port, 
      from_adder_to_mux_27_port, from_adder_to_mux_26_port, 
      from_adder_to_mux_25_port, from_adder_to_mux_24_port, 
      from_adder_to_mux_23_port, from_adder_to_mux_22_port, 
      from_adder_to_mux_21_port, from_adder_to_mux_20_port, 
      from_adder_to_mux_19_port, from_adder_to_mux_18_port, 
      from_adder_to_mux_17_port, from_adder_to_mux_16_port, 
      from_adder_to_mux_15_port, from_adder_to_mux_14_port, 
      from_adder_to_mux_13_port, from_adder_to_mux_12_port, 
      from_adder_to_mux_11_port, from_adder_to_mux_10_port, 
      from_adder_to_mux_9_port, from_adder_to_mux_8_port, 
      from_adder_to_mux_7_port, from_adder_to_mux_6_port, 
      from_adder_to_mux_5_port, from_adder_to_mux_4_port, 
      from_adder_to_mux_3_port, from_adder_to_mux_2_port, 
      from_adder_to_mux_1_port, from_adder_to_mux_0_port, 
      from_logict2_to_mux_31_port, from_logict2_to_mux_30_port, 
      from_logict2_to_mux_29_port, from_logict2_to_mux_28_port, 
      from_logict2_to_mux_27_port, from_logict2_to_mux_26_port, 
      from_logict2_to_mux_25_port, from_logict2_to_mux_24_port, 
      from_logict2_to_mux_23_port, from_logict2_to_mux_22_port, 
      from_logict2_to_mux_21_port, from_logict2_to_mux_20_port, 
      from_logict2_to_mux_19_port, from_logict2_to_mux_18_port, 
      from_logict2_to_mux_17_port, from_logict2_to_mux_16_port, 
      from_logict2_to_mux_15_port, from_logict2_to_mux_14_port, 
      from_logict2_to_mux_13_port, from_logict2_to_mux_12_port, 
      from_logict2_to_mux_11_port, from_logict2_to_mux_10_port, 
      from_logict2_to_mux_9_port, from_logict2_to_mux_8_port, 
      from_logict2_to_mux_7_port, from_logict2_to_mux_6_port, 
      from_logict2_to_mux_5_port, from_logict2_to_mux_4_port, 
      from_logict2_to_mux_3_port, from_logict2_to_mux_2_port, 
      from_logict2_to_mux_1_port, from_logict2_to_mux_0_port, 
      from_comparator_to_mux_31_port, from_comparator_to_mux_30_port, 
      from_comparator_to_mux_29_port, from_comparator_to_mux_28_port, 
      from_comparator_to_mux_27_port, from_comparator_to_mux_26_port, 
      from_comparator_to_mux_25_port, from_comparator_to_mux_24_port, 
      from_comparator_to_mux_23_port, from_comparator_to_mux_22_port, 
      from_comparator_to_mux_21_port, from_comparator_to_mux_20_port, 
      from_comparator_to_mux_19_port, from_comparator_to_mux_18_port, 
      from_comparator_to_mux_17_port, from_comparator_to_mux_16_port, 
      from_comparator_to_mux_15_port, from_comparator_to_mux_14_port, 
      from_comparator_to_mux_13_port, from_comparator_to_mux_12_port, 
      from_comparator_to_mux_11_port, from_comparator_to_mux_10_port, 
      from_comparator_to_mux_9_port, from_comparator_to_mux_8_port, 
      from_comparator_to_mux_7_port, from_comparator_to_mux_6_port, 
      from_comparator_to_mux_5_port, from_comparator_to_mux_4_port, 
      from_comparator_to_mux_3_port, from_comparator_to_mux_2_port, 
      from_comparator_to_mux_1_port, from_latch_to_logict2_op1_31_port, 
      from_latch_to_logict2_op1_30_port, from_latch_to_logict2_op1_29_port, 
      from_latch_to_logict2_op1_28_port, from_latch_to_logict2_op1_27_port, 
      from_latch_to_logict2_op1_26_port, from_latch_to_logict2_op1_25_port, 
      from_latch_to_logict2_op1_24_port, from_latch_to_logict2_op1_23_port, 
      from_latch_to_logict2_op1_22_port, from_latch_to_logict2_op1_21_port, 
      from_latch_to_logict2_op1_20_port, from_latch_to_logict2_op1_19_port, 
      from_latch_to_logict2_op1_18_port, from_latch_to_logict2_op1_17_port, 
      from_latch_to_logict2_op1_16_port, from_latch_to_logict2_op1_15_port, 
      from_latch_to_logict2_op1_14_port, from_latch_to_logict2_op1_13_port, 
      from_latch_to_logict2_op1_12_port, from_latch_to_logict2_op1_11_port, 
      from_latch_to_logict2_op1_10_port, from_latch_to_logict2_op1_9_port, 
      from_latch_to_logict2_op1_8_port, from_latch_to_logict2_op1_7_port, 
      from_latch_to_logict2_op1_6_port, from_latch_to_logict2_op1_5_port, 
      from_latch_to_logict2_op1_4_port, from_latch_to_logict2_op1_3_port, 
      from_latch_to_logict2_op1_2_port, from_latch_to_logict2_op1_1_port, 
      from_latch_to_logict2_op1_0_port, from_latch_to_logict2_op2_31_port, 
      from_latch_to_logict2_op2_30_port, from_latch_to_logict2_op2_29_port, 
      from_latch_to_logict2_op2_28_port, from_latch_to_logict2_op2_27_port, 
      from_latch_to_logict2_op2_26_port, from_latch_to_logict2_op2_25_port, 
      from_latch_to_logict2_op2_24_port, from_latch_to_logict2_op2_23_port, 
      from_latch_to_logict2_op2_22_port, from_latch_to_logict2_op2_21_port, 
      from_latch_to_logict2_op2_20_port, from_latch_to_logict2_op2_19_port, 
      from_latch_to_logict2_op2_18_port, from_latch_to_logict2_op2_17_port, 
      from_latch_to_logict2_op2_16_port, from_latch_to_logict2_op2_15_port, 
      from_latch_to_logict2_op2_14_port, from_latch_to_logict2_op2_13_port, 
      from_latch_to_logict2_op2_12_port, from_latch_to_logict2_op2_11_port, 
      from_latch_to_logict2_op2_10_port, from_latch_to_logict2_op2_9_port, 
      from_latch_to_logict2_op2_8_port, from_latch_to_logict2_op2_7_port, 
      from_latch_to_logict2_op2_6_port, from_latch_to_logict2_op2_5_port, 
      from_latch_to_logict2_op2_4_port, from_latch_to_logict2_op2_3_port, 
      from_latch_to_logict2_op2_2_port, from_latch_to_logict2_op2_1_port, 
      from_latch_to_logict2_op2_0_port, from_latch_to_comparator_op1_31_port, 
      from_latch_to_comparator_op1_30_port, 
      from_latch_to_comparator_op1_29_port, 
      from_latch_to_comparator_op1_28_port, 
      from_latch_to_comparator_op1_27_port, 
      from_latch_to_comparator_op1_26_port, 
      from_latch_to_comparator_op1_25_port, 
      from_latch_to_comparator_op1_24_port, 
      from_latch_to_comparator_op1_23_port, 
      from_latch_to_comparator_op1_22_port, 
      from_latch_to_comparator_op1_21_port, 
      from_latch_to_comparator_op1_20_port, 
      from_latch_to_comparator_op1_19_port, 
      from_latch_to_comparator_op1_18_port, 
      from_latch_to_comparator_op1_17_port, 
      from_latch_to_comparator_op1_16_port, 
      from_latch_to_comparator_op1_15_port, 
      from_latch_to_comparator_op1_14_port, 
      from_latch_to_comparator_op1_13_port, 
      from_latch_to_comparator_op1_12_port, 
      from_latch_to_comparator_op1_11_port, 
      from_latch_to_comparator_op1_10_port, from_latch_to_comparator_op1_9_port
      , from_latch_to_comparator_op1_8_port, 
      from_latch_to_comparator_op1_7_port, from_latch_to_comparator_op1_6_port,
      from_latch_to_comparator_op1_5_port, from_latch_to_comparator_op1_4_port,
      from_latch_to_comparator_op1_3_port, from_latch_to_comparator_op1_2_port,
      from_latch_to_comparator_op1_1_port, from_latch_to_comparator_op1_0_port,
      from_latch_to_comparator_op2_31_port, 
      from_latch_to_comparator_op2_30_port, 
      from_latch_to_comparator_op2_29_port, 
      from_latch_to_comparator_op2_28_port, 
      from_latch_to_comparator_op2_27_port, 
      from_latch_to_comparator_op2_26_port, 
      from_latch_to_comparator_op2_25_port, 
      from_latch_to_comparator_op2_24_port, 
      from_latch_to_comparator_op2_23_port, 
      from_latch_to_comparator_op2_22_port, 
      from_latch_to_comparator_op2_21_port, 
      from_latch_to_comparator_op2_20_port, 
      from_latch_to_comparator_op2_19_port, 
      from_latch_to_comparator_op2_18_port, 
      from_latch_to_comparator_op2_17_port, 
      from_latch_to_comparator_op2_16_port, 
      from_latch_to_comparator_op2_15_port, 
      from_latch_to_comparator_op2_14_port, 
      from_latch_to_comparator_op2_13_port, 
      from_latch_to_comparator_op2_12_port, 
      from_latch_to_comparator_op2_11_port, 
      from_latch_to_comparator_op2_10_port, from_latch_to_comparator_op2_9_port
      , from_latch_to_comparator_op2_8_port, 
      from_latch_to_comparator_op2_7_port, from_latch_to_comparator_op2_6_port,
      from_latch_to_comparator_op2_5_port, from_latch_to_comparator_op2_4_port,
      from_latch_to_comparator_op2_3_port, from_latch_to_comparator_op2_2_port,
      from_latch_to_comparator_op2_1_port, from_latch_to_comparator_op2_0_port,
      net2772, net2773, net2774, net2775, net2776, net2777, net2778, net2779, 
      net2780, net2781, net2782, net2783, net2784, net2785, net2786, net2787, 
      net2788, net2789, net2790, net2791, net2792, net2793, net2794, net2795, 
      net2796, net2797, net2798, net2799, net2800, net2801, net2802, net2803, 
      net2771, net2770, net2769, net2768, net2767, net2766, net2765, net2764, 
      net2763, net2762, net2761, net2760, net2759, net2758, net2757, net2756, 
      net2755, net2754, net2753, net2752, net2751, net2750, net2749, net2748, 
      net2747, net2746, net2745, net2744, net2743, net2742, net2741, net2740, 
      net2739, net2738, mux_to_mux_low_9_port, mux_to_mux_low_8_port, 
      mux_to_mux_low_7_port, mux_to_mux_low_6_port, mux_to_mux_low_5_port, 
      mux_to_mux_low_4_port, mux_to_mux_low_3_port, mux_to_mux_low_31_port, 
      mux_to_mux_low_30_port, mux_to_mux_low_2_port, mux_to_mux_low_29_port, 
      mux_to_mux_low_28_port, mux_to_mux_low_27_port, mux_to_mux_low_26_port, 
      mux_to_mux_low_25_port, mux_to_mux_low_24_port, mux_to_mux_low_23_port, 
      mux_to_mux_low_22_port, mux_to_mux_low_21_port, mux_to_mux_low_20_port, 
      mux_to_mux_low_1_port, mux_to_mux_low_19_port, mux_to_mux_low_18_port, 
      mux_to_mux_low_17_port, mux_to_mux_low_16_port, mux_to_mux_low_15_port, 
      mux_to_mux_low_14_port, mux_to_mux_low_13_port, mux_to_mux_low_12_port, 
      mux_to_mux_low_11_port, mux_to_mux_low_10_port, mux_to_mux_low_0_port, 
      mux_to_mux_high_9_port, mux_to_mux_high_8_port, mux_to_mux_high_7_port, 
      mux_to_mux_high_6_port, mux_to_mux_high_5_port, mux_to_mux_high_4_port, 
      mux_to_mux_high_3_port, mux_to_mux_high_31_port, mux_to_mux_high_30_port,
      mux_to_mux_high_2_port, mux_to_mux_high_29_port, mux_to_mux_high_28_port,
      mux_to_mux_high_27_port, mux_to_mux_high_26_port, mux_to_mux_high_25_port
      , mux_to_mux_high_24_port, mux_to_mux_high_23_port, 
      mux_to_mux_high_22_port, mux_to_mux_high_21_port, mux_to_mux_high_20_port
      , mux_to_mux_high_1_port, mux_to_mux_high_19_port, 
      mux_to_mux_high_18_port, mux_to_mux_high_17_port, mux_to_mux_high_16_port
      , mux_to_mux_high_15_port, mux_to_mux_high_14_port, 
      mux_to_mux_high_13_port, mux_to_mux_high_12_port, mux_to_mux_high_11_port
      , mux_to_mux_high_10_port, mux_to_mux_high_0_port, 
      from_mux_2_1_to_reg_9_port, from_mux_2_1_to_reg_8_port, 
      from_mux_2_1_to_reg_7_port, from_mux_2_1_to_reg_6_port, 
      from_mux_2_1_to_reg_5_port, from_mux_2_1_to_reg_4_port, 
      from_mux_2_1_to_reg_3_port, from_mux_2_1_to_reg_31_port, 
      from_mux_2_1_to_reg_30_port, from_mux_2_1_to_reg_2_port, 
      from_mux_2_1_to_reg_29_port, from_mux_2_1_to_reg_28_port, 
      from_mux_2_1_to_reg_27_port, from_mux_2_1_to_reg_26_port, 
      from_mux_2_1_to_reg_25_port, from_mux_2_1_to_reg_24_port, 
      from_mux_2_1_to_reg_23_port, from_mux_2_1_to_reg_22_port, 
      from_mux_2_1_to_reg_21_port, from_mux_2_1_to_reg_20_port, 
      from_mux_2_1_to_reg_1_port, from_mux_2_1_to_reg_19_port, 
      from_mux_2_1_to_reg_18_port, from_mux_2_1_to_reg_17_port, 
      from_mux_2_1_to_reg_16_port, from_mux_2_1_to_reg_15_port, 
      from_mux_2_1_to_reg_14_port, from_mux_2_1_to_reg_13_port, 
      from_mux_2_1_to_reg_12_port, from_mux_2_1_to_reg_11_port, 
      from_mux_2_1_to_reg_10_port, from_mux_2_1_to_reg_0_port, 
      from_latch_to_mux_sub_or_add_9_port, from_latch_to_mux_sub_or_add_8_port,
      from_latch_to_mux_sub_or_add_7_port, from_latch_to_mux_sub_or_add_6_port,
      from_latch_to_mux_sub_or_add_5_port, from_latch_to_mux_sub_or_add_4_port,
      from_latch_to_mux_sub_or_add_3_port, from_latch_to_mux_sub_or_add_31_port
      , from_latch_to_mux_sub_or_add_30_port, 
      from_latch_to_mux_sub_or_add_2_port, from_latch_to_mux_sub_or_add_29_port
      , from_latch_to_mux_sub_or_add_28_port, 
      from_latch_to_mux_sub_or_add_27_port, 
      from_latch_to_mux_sub_or_add_26_port, 
      from_latch_to_mux_sub_or_add_25_port, 
      from_latch_to_mux_sub_or_add_24_port, 
      from_latch_to_mux_sub_or_add_23_port, 
      from_latch_to_mux_sub_or_add_22_port, 
      from_latch_to_mux_sub_or_add_21_port, 
      from_latch_to_mux_sub_or_add_20_port, from_latch_to_mux_sub_or_add_1_port
      , from_latch_to_mux_sub_or_add_19_port, 
      from_latch_to_mux_sub_or_add_18_port, 
      from_latch_to_mux_sub_or_add_17_port, 
      from_latch_to_mux_sub_or_add_16_port, 
      from_latch_to_mux_sub_or_add_15_port, 
      from_latch_to_mux_sub_or_add_14_port, 
      from_latch_to_mux_sub_or_add_13_port, 
      from_latch_to_mux_sub_or_add_12_port, 
      from_latch_to_mux_sub_or_add_11_port, 
      from_latch_to_mux_sub_or_add_10_port, from_latch_to_mux_sub_or_add_0_port
      , from_latch_to_adder_op1_9_port, from_latch_to_adder_op1_8_port, 
      from_latch_to_adder_op1_7_port, from_latch_to_adder_op1_6_port, 
      from_latch_to_adder_op1_5_port, from_latch_to_adder_op1_4_port, 
      from_latch_to_adder_op1_3_port, from_latch_to_adder_op1_31_port, 
      from_latch_to_adder_op1_30_port, from_latch_to_adder_op1_2_port, 
      from_latch_to_adder_op1_29_port, from_latch_to_adder_op1_28_port, 
      from_latch_to_adder_op1_27_port, from_latch_to_adder_op1_26_port, 
      from_latch_to_adder_op1_25_port, from_latch_to_adder_op1_24_port, 
      from_latch_to_adder_op1_23_port, from_latch_to_adder_op1_22_port, 
      from_latch_to_adder_op1_21_port, from_latch_to_adder_op1_20_port, 
      from_latch_to_adder_op1_1_port, from_latch_to_adder_op1_19_port, 
      from_latch_to_adder_op1_18_port, from_latch_to_adder_op1_17_port, 
      from_latch_to_adder_op1_16_port, from_latch_to_adder_op1_15_port, 
      from_latch_to_adder_op1_14_port, from_latch_to_adder_op1_13_port, 
      from_latch_to_adder_op1_12_port, from_latch_to_adder_op1_11_port, 
      from_latch_to_adder_op1_10_port, from_latch_to_adder_op1_0_port, n4, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086 : std_logic;

begin
   jump <= jump_port;
   
   from_comparator_to_mux_1_port <= '0';
   from_comparator_to_mux_2_port <= '0';
   from_comparator_to_mux_3_port <= '0';
   from_comparator_to_mux_4_port <= '0';
   from_comparator_to_mux_5_port <= '0';
   from_comparator_to_mux_6_port <= '0';
   from_comparator_to_mux_7_port <= '0';
   from_comparator_to_mux_8_port <= '0';
   from_comparator_to_mux_9_port <= '0';
   from_comparator_to_mux_10_port <= '0';
   from_comparator_to_mux_11_port <= '0';
   from_comparator_to_mux_12_port <= '0';
   from_comparator_to_mux_13_port <= '0';
   from_comparator_to_mux_14_port <= '0';
   from_comparator_to_mux_15_port <= '0';
   from_comparator_to_mux_16_port <= '0';
   from_comparator_to_mux_17_port <= '0';
   from_comparator_to_mux_18_port <= '0';
   from_comparator_to_mux_19_port <= '0';
   from_comparator_to_mux_20_port <= '0';
   from_comparator_to_mux_21_port <= '0';
   from_comparator_to_mux_22_port <= '0';
   from_comparator_to_mux_23_port <= '0';
   from_comparator_to_mux_24_port <= '0';
   from_comparator_to_mux_25_port <= '0';
   from_comparator_to_mux_26_port <= '0';
   from_comparator_to_mux_27_port <= '0';
   from_comparator_to_mux_28_port <= '0';
   from_comparator_to_mux_29_port <= '0';
   from_comparator_to_mux_30_port <= '0';
   from_comparator_to_mux_31_port <= '0';
   signal_cmd_t2_0_port <= '0';
   RE_2 : regWithEnable_6 port map( input(31) => mux_to_mux_low_31_port, 
                           input(30) => mux_to_mux_low_30_port, input(29) => 
                           mux_to_mux_low_29_port, input(28) => 
                           mux_to_mux_low_28_port, input(27) => 
                           mux_to_mux_low_27_port, input(26) => 
                           mux_to_mux_low_26_port, input(25) => 
                           mux_to_mux_low_25_port, input(24) => 
                           mux_to_mux_low_24_port, input(23) => 
                           mux_to_mux_low_23_port, input(22) => 
                           mux_to_mux_low_22_port, input(21) => 
                           mux_to_mux_low_21_port, input(20) => 
                           mux_to_mux_low_20_port, input(19) => 
                           mux_to_mux_low_19_port, input(18) => 
                           mux_to_mux_low_18_port, input(17) => 
                           mux_to_mux_low_17_port, input(16) => 
                           mux_to_mux_low_16_port, input(15) => 
                           mux_to_mux_low_15_port, input(14) => 
                           mux_to_mux_low_14_port, input(13) => 
                           mux_to_mux_low_13_port, input(12) => 
                           mux_to_mux_low_12_port, input(11) => 
                           mux_to_mux_low_11_port, input(10) => 
                           mux_to_mux_low_10_port, input(9) => 
                           mux_to_mux_low_9_port, input(8) => 
                           mux_to_mux_low_8_port, input(7) => 
                           mux_to_mux_low_7_port, input(6) => 
                           mux_to_mux_low_6_port, input(5) => 
                           mux_to_mux_low_5_port, input(4) => 
                           mux_to_mux_low_4_port, input(3) => 
                           mux_to_mux_low_3_port, input(2) => 
                           mux_to_mux_low_2_port, input(1) => 
                           mux_to_mux_low_1_port, input(0) => 
                           mux_to_mux_low_0_port, en => enable, clock => clock,
                           reset => reset, output(31) => 
                           out_res_operand_two(31), output(30) => 
                           out_res_operand_two(30), output(29) => 
                           out_res_operand_two(29), output(28) => 
                           out_res_operand_two(28), output(27) => 
                           out_res_operand_two(27), output(26) => 
                           out_res_operand_two(26), output(25) => 
                           out_res_operand_two(25), output(24) => 
                           out_res_operand_two(24), output(23) => 
                           out_res_operand_two(23), output(22) => 
                           out_res_operand_two(22), output(21) => 
                           out_res_operand_two(21), output(20) => 
                           out_res_operand_two(20), output(19) => 
                           out_res_operand_two(19), output(18) => 
                           out_res_operand_two(18), output(17) => 
                           out_res_operand_two(17), output(16) => 
                           out_res_operand_two(16), output(15) => 
                           out_res_operand_two(15), output(14) => 
                           out_res_operand_two(14), output(13) => 
                           out_res_operand_two(13), output(12) => 
                           out_res_operand_two(12), output(11) => 
                           out_res_operand_two(11), output(10) => 
                           out_res_operand_two(10), output(9) => 
                           out_res_operand_two(9), output(8) => 
                           out_res_operand_two(8), output(7) => 
                           out_res_operand_two(7), output(6) => 
                           out_res_operand_two(6), output(5) => 
                           out_res_operand_two(5), output(4) => 
                           out_res_operand_two(4), output(3) => 
                           out_res_operand_two(3), output(2) => 
                           out_res_operand_two(2), output(1) => 
                           out_res_operand_two(1), output(0) => 
                           out_res_operand_two(0));
   CU_EX : cu_exe port map( reset => reset, func(10) => func(10), func(9) => 
                           func(9), func(8) => func(8), func(7) => func(7), 
                           func(6) => func(6), func(5) => func(5), func(4) => 
                           func(4), func(3) => func(3), func(2) => func(2), 
                           func(1) => func(1), func(0) => func(0), busy_div => 
                           busy, multi_cycle_operation => multi_cycle_operation
                           , enable => enable_mux_4_1, sel_signal_5X1(2) => 
                           sel_signal_5_1_2_port, sel_signal_5X1(1) => 
                           sel_signal_5_1_1_port, sel_signal_5X1(0) => 
                           sel_signal_5_1_0_port, sel_signal_2X1 => 
                           sel_signal_2_1, start_div => start_div, cmd_t2(3) =>
                           signal_cmd_t2_3_port, cmd_t2(2) => 
                           signal_cmd_t2_2_port, cmd_t2(1) => 
                           signal_cmd_t2_1_port, cmd_t2(0) => n_1055, carry_in 
                           => carry_in, left_right => left_right, logic_Arith 
                           => logic_Arith, shift_rot => shift_rot, 
                           sel_comparator(2) => sel_comparator_2_port, 
                           sel_comparator(1) => sel_comparator_1_port, 
                           sel_comparator(0) => sel_comparator_0_port);
   RE_1 : regWithEnable_5bit_4 port map( input(4) => EX_MEM_rd_next_4_port, 
                           input(3) => EX_MEM_rd_next_3_port, input(2) => 
                           EX_MEM_rd_next_2_port, input(1) => 
                           EX_MEM_rd_next_1_port, input(0) => 
                           EX_MEM_rd_next_0_port, en => enable, clock => clock,
                           reset => reset, output(4) => EX_MEM_rd(4), output(3)
                           => EX_MEM_rd(3), output(2) => EX_MEM_rd(2), 
                           output(1) => EX_MEM_rd(1), output(0) => EX_MEM_rd(0)
                           );
   M6 : mux_2_1_5bit port map( a(4) => ID_EX_Rd(4), a(3) => ID_EX_Rd(3), a(2) 
                           => ID_EX_Rd(2), a(1) => ID_EX_Rd(1), a(0) => 
                           ID_EX_Rd(0), b(4) => ID_EX_Rt(4), b(3) => 
                           ID_EX_Rt(3), b(2) => ID_EX_Rt(2), b(1) => 
                           ID_EX_Rt(1), b(0) => ID_EX_Rt(0), sel => sel_3, o(4)
                           => EX_MEM_rd_next_4_port, o(3) => 
                           EX_MEM_rd_next_3_port, o(2) => EX_MEM_rd_next_2_port
                           , o(1) => EX_MEM_rd_next_1_port, o(0) => 
                           EX_MEM_rd_next_0_port);
   FU : forwarding_unit port map( EX_MEM_write => EX_MEM_write, EX_MEM_Rd(4) =>
                           EX_MEM_rd(4), EX_MEM_Rd(3) => EX_MEM_rd(3), 
                           EX_MEM_Rd(2) => EX_MEM_rd(2), EX_MEM_Rd(1) => 
                           EX_MEM_rd(1), EX_MEM_Rd(0) => EX_MEM_rd(0), 
                           ID_EX_Rs(4) => ID_EX_Rs(4), ID_EX_Rs(3) => 
                           ID_EX_Rs(3), ID_EX_Rs(2) => ID_EX_Rs(2), ID_EX_Rs(1)
                           => ID_EX_Rs(1), ID_EX_Rs(0) => ID_EX_Rs(0), 
                           ID_EX_Rt(4) => ID_EX_Rt(4), ID_EX_Rt(3) => 
                           ID_EX_Rt(3), ID_EX_Rt(2) => ID_EX_Rt(2), ID_EX_Rt(1)
                           => ID_EX_Rt(1), ID_EX_Rt(0) => ID_EX_Rt(0), 
                           MEM_WB_write => MEM_WB_write, MEM_WB_Rd(4) => 
                           MEM_WB_rd(4), MEM_WB_Rd(3) => MEM_WB_rd(3), 
                           MEM_WB_Rd(2) => MEM_WB_rd(2), MEM_WB_Rd(1) => 
                           MEM_WB_rd(1), MEM_WB_Rd(0) => MEM_WB_rd(0), 
                           sel_mux_high(1) => sel_mux_3_1_high_1_port, 
                           sel_mux_high(0) => sel_mux_3_1_high_0_port, 
                           sel_mux_low(1) => sel_mux_3_1_low_1_port, 
                           sel_mux_low(0) => sel_mux_3_1_low_0_port);
   M5 : Mux2X1_5 port map( a(31) => quotient_31_port, a(30) => quotient_30_port
                           , a(29) => quotient_29_port, a(28) => 
                           quotient_28_port, a(27) => quotient_27_port, a(26) 
                           => quotient_26_port, a(25) => quotient_25_port, 
                           a(24) => quotient_24_port, a(23) => quotient_23_port
                           , a(22) => quotient_22_port, a(21) => 
                           quotient_21_port, a(20) => quotient_20_port, a(19) 
                           => quotient_19_port, a(18) => quotient_18_port, 
                           a(17) => quotient_17_port, a(16) => quotient_16_port
                           , a(15) => quotient_15_port, a(14) => 
                           quotient_14_port, a(13) => quotient_13_port, a(12) 
                           => quotient_12_port, a(11) => quotient_11_port, 
                           a(10) => quotient_10_port, a(9) => quotient_9_port, 
                           a(8) => quotient_8_port, a(7) => quotient_7_port, 
                           a(6) => quotient_6_port, a(5) => quotient_5_port, 
                           a(4) => quotient_4_port, a(3) => quotient_3_port, 
                           a(2) => quotient_2_port, a(1) => quotient_1_port, 
                           a(0) => quotient_0_port, b(31) => 
                           from_mux_4_1_to_mux_2_1_31_port, b(30) => 
                           from_mux_4_1_to_mux_2_1_30_port, b(29) => 
                           from_mux_4_1_to_mux_2_1_29_port, b(28) => 
                           from_mux_4_1_to_mux_2_1_28_port, b(27) => 
                           from_mux_4_1_to_mux_2_1_27_port, b(26) => 
                           from_mux_4_1_to_mux_2_1_26_port, b(25) => 
                           from_mux_4_1_to_mux_2_1_25_port, b(24) => 
                           from_mux_4_1_to_mux_2_1_24_port, b(23) => 
                           from_mux_4_1_to_mux_2_1_23_port, b(22) => 
                           from_mux_4_1_to_mux_2_1_22_port, b(21) => 
                           from_mux_4_1_to_mux_2_1_21_port, b(20) => 
                           from_mux_4_1_to_mux_2_1_20_port, b(19) => 
                           from_mux_4_1_to_mux_2_1_19_port, b(18) => 
                           from_mux_4_1_to_mux_2_1_18_port, b(17) => 
                           from_mux_4_1_to_mux_2_1_17_port, b(16) => 
                           from_mux_4_1_to_mux_2_1_16_port, b(15) => 
                           from_mux_4_1_to_mux_2_1_15_port, b(14) => 
                           from_mux_4_1_to_mux_2_1_14_port, b(13) => 
                           from_mux_4_1_to_mux_2_1_13_port, b(12) => 
                           from_mux_4_1_to_mux_2_1_12_port, b(11) => 
                           from_mux_4_1_to_mux_2_1_11_port, b(10) => 
                           from_mux_4_1_to_mux_2_1_10_port, b(9) => 
                           from_mux_4_1_to_mux_2_1_9_port, b(8) => 
                           from_mux_4_1_to_mux_2_1_8_port, b(7) => 
                           from_mux_4_1_to_mux_2_1_7_port, b(6) => 
                           from_mux_4_1_to_mux_2_1_6_port, b(5) => 
                           from_mux_4_1_to_mux_2_1_5_port, b(4) => 
                           from_mux_4_1_to_mux_2_1_4_port, b(3) => 
                           from_mux_4_1_to_mux_2_1_3_port, b(2) => 
                           from_mux_4_1_to_mux_2_1_2_port, b(1) => 
                           from_mux_4_1_to_mux_2_1_1_port, b(0) => 
                           from_mux_4_1_to_mux_2_1_0_port, sel => 
                           sel_signal_2_1, o(31) => from_mux_2_1_to_reg_31_port
                           , o(30) => from_mux_2_1_to_reg_30_port, o(29) => 
                           from_mux_2_1_to_reg_29_port, o(28) => 
                           from_mux_2_1_to_reg_28_port, o(27) => 
                           from_mux_2_1_to_reg_27_port, o(26) => 
                           from_mux_2_1_to_reg_26_port, o(25) => 
                           from_mux_2_1_to_reg_25_port, o(24) => 
                           from_mux_2_1_to_reg_24_port, o(23) => 
                           from_mux_2_1_to_reg_23_port, o(22) => 
                           from_mux_2_1_to_reg_22_port, o(21) => 
                           from_mux_2_1_to_reg_21_port, o(20) => 
                           from_mux_2_1_to_reg_20_port, o(19) => 
                           from_mux_2_1_to_reg_19_port, o(18) => 
                           from_mux_2_1_to_reg_18_port, o(17) => 
                           from_mux_2_1_to_reg_17_port, o(16) => 
                           from_mux_2_1_to_reg_16_port, o(15) => 
                           from_mux_2_1_to_reg_15_port, o(14) => 
                           from_mux_2_1_to_reg_14_port, o(13) => 
                           from_mux_2_1_to_reg_13_port, o(12) => 
                           from_mux_2_1_to_reg_12_port, o(11) => 
                           from_mux_2_1_to_reg_11_port, o(10) => 
                           from_mux_2_1_to_reg_10_port, o(9) => 
                           from_mux_2_1_to_reg_9_port, o(8) => 
                           from_mux_2_1_to_reg_8_port, o(7) => 
                           from_mux_2_1_to_reg_7_port, o(6) => 
                           from_mux_2_1_to_reg_6_port, o(5) => 
                           from_mux_2_1_to_reg_5_port, o(4) => 
                           from_mux_2_1_to_reg_4_port, o(3) => 
                           from_mux_2_1_to_reg_3_port, o(2) => 
                           from_mux_2_1_to_reg_2_port, o(1) => 
                           from_mux_2_1_to_reg_1_port, o(0) => 
                           from_mux_2_1_to_reg_0_port);
   DM : DIVIDER_N_op32 port map( CLK => clock, START => start_div, RESET => 
                           reset, BUSY => busy, DIVIDEND(31) => 
                           from_mux_2_1_to_latch_high_31_port, DIVIDEND(30) => 
                           from_mux_2_1_to_latch_high_30_port, DIVIDEND(29) => 
                           from_mux_2_1_to_latch_high_29_port, DIVIDEND(28) => 
                           from_mux_2_1_to_latch_high_28_port, DIVIDEND(27) => 
                           from_mux_2_1_to_latch_high_27_port, DIVIDEND(26) => 
                           from_mux_2_1_to_latch_high_26_port, DIVIDEND(25) => 
                           from_mux_2_1_to_latch_high_25_port, DIVIDEND(24) => 
                           from_mux_2_1_to_latch_high_24_port, DIVIDEND(23) => 
                           from_mux_2_1_to_latch_high_23_port, DIVIDEND(22) => 
                           from_mux_2_1_to_latch_high_22_port, DIVIDEND(21) => 
                           from_mux_2_1_to_latch_high_21_port, DIVIDEND(20) => 
                           from_mux_2_1_to_latch_high_20_port, DIVIDEND(19) => 
                           from_mux_2_1_to_latch_high_19_port, DIVIDEND(18) => 
                           from_mux_2_1_to_latch_high_18_port, DIVIDEND(17) => 
                           from_mux_2_1_to_latch_high_17_port, DIVIDEND(16) => 
                           from_mux_2_1_to_latch_high_16_port, DIVIDEND(15) => 
                           from_mux_2_1_to_latch_high_15_port, DIVIDEND(14) => 
                           from_mux_2_1_to_latch_high_14_port, DIVIDEND(13) => 
                           from_mux_2_1_to_latch_high_13_port, DIVIDEND(12) => 
                           from_mux_2_1_to_latch_high_12_port, DIVIDEND(11) => 
                           from_mux_2_1_to_latch_high_11_port, DIVIDEND(10) => 
                           from_mux_2_1_to_latch_high_10_port, DIVIDEND(9) => 
                           from_mux_2_1_to_latch_high_9_port, DIVIDEND(8) => 
                           from_mux_2_1_to_latch_high_8_port, DIVIDEND(7) => 
                           from_mux_2_1_to_latch_high_7_port, DIVIDEND(6) => 
                           from_mux_2_1_to_latch_high_6_port, DIVIDEND(5) => 
                           from_mux_2_1_to_latch_high_5_port, DIVIDEND(4) => 
                           from_mux_2_1_to_latch_high_4_port, DIVIDEND(3) => 
                           from_mux_2_1_to_latch_high_3_port, DIVIDEND(2) => 
                           from_mux_2_1_to_latch_high_2_port, DIVIDEND(1) => 
                           from_mux_2_1_to_latch_high_1_port, DIVIDEND(0) => 
                           from_mux_2_1_to_latch_high_0_port, DIVISOR(31) => 
                           from_mux_2_1_to_latch_low_31_port, DIVISOR(30) => 
                           from_mux_2_1_to_latch_low_30_port, DIVISOR(29) => 
                           from_mux_2_1_to_latch_low_29_port, DIVISOR(28) => 
                           from_mux_2_1_to_latch_low_28_port, DIVISOR(27) => 
                           from_mux_2_1_to_latch_low_27_port, DIVISOR(26) => 
                           from_mux_2_1_to_latch_low_26_port, DIVISOR(25) => 
                           from_mux_2_1_to_latch_low_25_port, DIVISOR(24) => 
                           from_mux_2_1_to_latch_low_24_port, DIVISOR(23) => 
                           from_mux_2_1_to_latch_low_23_port, DIVISOR(22) => 
                           from_mux_2_1_to_latch_low_22_port, DIVISOR(21) => 
                           from_mux_2_1_to_latch_low_21_port, DIVISOR(20) => 
                           from_mux_2_1_to_latch_low_20_port, DIVISOR(19) => 
                           from_mux_2_1_to_latch_low_19_port, DIVISOR(18) => 
                           from_mux_2_1_to_latch_low_18_port, DIVISOR(17) => 
                           from_mux_2_1_to_latch_low_17_port, DIVISOR(16) => 
                           from_mux_2_1_to_latch_low_16_port, DIVISOR(15) => 
                           from_mux_2_1_to_latch_low_15_port, DIVISOR(14) => 
                           from_mux_2_1_to_latch_low_14_port, DIVISOR(13) => 
                           from_mux_2_1_to_latch_low_13_port, DIVISOR(12) => 
                           from_mux_2_1_to_latch_low_12_port, DIVISOR(11) => 
                           from_mux_2_1_to_latch_low_11_port, DIVISOR(10) => 
                           from_mux_2_1_to_latch_low_10_port, DIVISOR(9) => 
                           from_mux_2_1_to_latch_low_9_port, DIVISOR(8) => 
                           from_mux_2_1_to_latch_low_8_port, DIVISOR(7) => 
                           from_mux_2_1_to_latch_low_7_port, DIVISOR(6) => 
                           from_mux_2_1_to_latch_low_6_port, DIVISOR(5) => 
                           from_mux_2_1_to_latch_low_5_port, DIVISOR(4) => 
                           from_mux_2_1_to_latch_low_4_port, DIVISOR(3) => 
                           from_mux_2_1_to_latch_low_3_port, DIVISOR(2) => 
                           from_mux_2_1_to_latch_low_2_port, DIVISOR(1) => 
                           from_mux_2_1_to_latch_low_1_port, DIVISOR(0) => 
                           from_mux_2_1_to_latch_low_0_port, QUOTIENT(31) => 
                           quotient_31_port, QUOTIENT(30) => quotient_30_port, 
                           QUOTIENT(29) => quotient_29_port, QUOTIENT(28) => 
                           quotient_28_port, QUOTIENT(27) => quotient_27_port, 
                           QUOTIENT(26) => quotient_26_port, QUOTIENT(25) => 
                           quotient_25_port, QUOTIENT(24) => quotient_24_port, 
                           QUOTIENT(23) => quotient_23_port, QUOTIENT(22) => 
                           quotient_22_port, QUOTIENT(21) => quotient_21_port, 
                           QUOTIENT(20) => quotient_20_port, QUOTIENT(19) => 
                           quotient_19_port, QUOTIENT(18) => quotient_18_port, 
                           QUOTIENT(17) => quotient_17_port, QUOTIENT(16) => 
                           quotient_16_port, QUOTIENT(15) => quotient_15_port, 
                           QUOTIENT(14) => quotient_14_port, QUOTIENT(13) => 
                           quotient_13_port, QUOTIENT(12) => quotient_12_port, 
                           QUOTIENT(11) => quotient_11_port, QUOTIENT(10) => 
                           quotient_10_port, QUOTIENT(9) => quotient_9_port, 
                           QUOTIENT(8) => quotient_8_port, QUOTIENT(7) => 
                           quotient_7_port, QUOTIENT(6) => quotient_6_port, 
                           QUOTIENT(5) => quotient_5_port, QUOTIENT(4) => 
                           quotient_4_port, QUOTIENT(3) => quotient_3_port, 
                           QUOTIENT(2) => quotient_2_port, QUOTIENT(1) => 
                           quotient_1_port, QUOTIENT(0) => quotient_0_port, 
                           RESIDUAL(31) => net2772, RESIDUAL(30) => net2773, 
                           RESIDUAL(29) => net2774, RESIDUAL(28) => net2775, 
                           RESIDUAL(27) => net2776, RESIDUAL(26) => net2777, 
                           RESIDUAL(25) => net2778, RESIDUAL(24) => net2779, 
                           RESIDUAL(23) => net2780, RESIDUAL(22) => net2781, 
                           RESIDUAL(21) => net2782, RESIDUAL(20) => net2783, 
                           RESIDUAL(19) => net2784, RESIDUAL(18) => net2785, 
                           RESIDUAL(17) => net2786, RESIDUAL(16) => net2787, 
                           RESIDUAL(15) => net2788, RESIDUAL(14) => net2789, 
                           RESIDUAL(13) => net2790, RESIDUAL(12) => net2791, 
                           RESIDUAL(11) => net2792, RESIDUAL(10) => net2793, 
                           RESIDUAL(9) => net2794, RESIDUAL(8) => net2795, 
                           RESIDUAL(7) => net2796, RESIDUAL(6) => net2797, 
                           RESIDUAL(5) => net2798, RESIDUAL(4) => net2799, 
                           RESIDUAL(3) => net2800, RESIDUAL(2) => net2801, 
                           RESIDUAL(1) => net2802, RESIDUAL(0) => net2803);
   RE : regWithEnable_5 port map( input(31) => from_mux_2_1_to_reg_31_port, 
                           input(30) => from_mux_2_1_to_reg_30_port, input(29) 
                           => from_mux_2_1_to_reg_29_port, input(28) => 
                           from_mux_2_1_to_reg_28_port, input(27) => 
                           from_mux_2_1_to_reg_27_port, input(26) => 
                           from_mux_2_1_to_reg_26_port, input(25) => 
                           from_mux_2_1_to_reg_25_port, input(24) => 
                           from_mux_2_1_to_reg_24_port, input(23) => 
                           from_mux_2_1_to_reg_23_port, input(22) => 
                           from_mux_2_1_to_reg_22_port, input(21) => 
                           from_mux_2_1_to_reg_21_port, input(20) => 
                           from_mux_2_1_to_reg_20_port, input(19) => 
                           from_mux_2_1_to_reg_19_port, input(18) => 
                           from_mux_2_1_to_reg_18_port, input(17) => 
                           from_mux_2_1_to_reg_17_port, input(16) => 
                           from_mux_2_1_to_reg_16_port, input(15) => 
                           from_mux_2_1_to_reg_15_port, input(14) => 
                           from_mux_2_1_to_reg_14_port, input(13) => 
                           from_mux_2_1_to_reg_13_port, input(12) => 
                           from_mux_2_1_to_reg_12_port, input(11) => 
                           from_mux_2_1_to_reg_11_port, input(10) => 
                           from_mux_2_1_to_reg_10_port, input(9) => 
                           from_mux_2_1_to_reg_9_port, input(8) => 
                           from_mux_2_1_to_reg_8_port, input(7) => 
                           from_mux_2_1_to_reg_7_port, input(6) => 
                           from_mux_2_1_to_reg_6_port, input(5) => 
                           from_mux_2_1_to_reg_5_port, input(4) => 
                           from_mux_2_1_to_reg_4_port, input(3) => 
                           from_mux_2_1_to_reg_3_port, input(2) => 
                           from_mux_2_1_to_reg_2_port, input(1) => 
                           from_mux_2_1_to_reg_1_port, input(0) => 
                           from_mux_2_1_to_reg_0_port, en => enable, clock => 
                           clock, reset => reset, output(31) => 
                           out_res_operand_one(31), output(30) => 
                           out_res_operand_one(30), output(29) => 
                           out_res_operand_one(29), output(28) => 
                           out_res_operand_one(28), output(27) => 
                           out_res_operand_one(27), output(26) => 
                           out_res_operand_one(26), output(25) => 
                           out_res_operand_one(25), output(24) => 
                           out_res_operand_one(24), output(23) => 
                           out_res_operand_one(23), output(22) => 
                           out_res_operand_one(22), output(21) => 
                           out_res_operand_one(21), output(20) => 
                           out_res_operand_one(20), output(19) => 
                           out_res_operand_one(19), output(18) => 
                           out_res_operand_one(18), output(17) => 
                           out_res_operand_one(17), output(16) => 
                           out_res_operand_one(16), output(15) => 
                           out_res_operand_one(15), output(14) => 
                           out_res_operand_one(14), output(13) => 
                           out_res_operand_one(13), output(12) => 
                           out_res_operand_one(12), output(11) => 
                           out_res_operand_one(11), output(10) => 
                           out_res_operand_one(10), output(9) => 
                           out_res_operand_one(9), output(8) => 
                           out_res_operand_one(8), output(7) => 
                           out_res_operand_one(7), output(6) => 
                           out_res_operand_one(6), output(5) => 
                           out_res_operand_one(5), output(4) => 
                           out_res_operand_one(4), output(3) => 
                           out_res_operand_one(3), output(2) => 
                           out_res_operand_one(2), output(1) => 
                           out_res_operand_one(1), output(0) => 
                           out_res_operand_one(0));
   SF : Shifter_NBIT32 port map( left_right => left_right, logic_Arith => 
                           logic_Arith, shift_rot => shift_rot, a(31) => 
                           from_latch_to_shifter_op1_31_port, a(30) => 
                           from_latch_to_shifter_op1_30_port, a(29) => 
                           from_latch_to_shifter_op1_29_port, a(28) => 
                           from_latch_to_shifter_op1_28_port, a(27) => 
                           from_latch_to_shifter_op1_27_port, a(26) => 
                           from_latch_to_shifter_op1_26_port, a(25) => 
                           from_latch_to_shifter_op1_25_port, a(24) => 
                           from_latch_to_shifter_op1_24_port, a(23) => 
                           from_latch_to_shifter_op1_23_port, a(22) => 
                           from_latch_to_shifter_op1_22_port, a(21) => 
                           from_latch_to_shifter_op1_21_port, a(20) => 
                           from_latch_to_shifter_op1_20_port, a(19) => 
                           from_latch_to_shifter_op1_19_port, a(18) => 
                           from_latch_to_shifter_op1_18_port, a(17) => 
                           from_latch_to_shifter_op1_17_port, a(16) => 
                           from_latch_to_shifter_op1_16_port, a(15) => 
                           from_latch_to_shifter_op1_15_port, a(14) => 
                           from_latch_to_shifter_op1_14_port, a(13) => 
                           from_latch_to_shifter_op1_13_port, a(12) => 
                           from_latch_to_shifter_op1_12_port, a(11) => 
                           from_latch_to_shifter_op1_11_port, a(10) => 
                           from_latch_to_shifter_op1_10_port, a(9) => 
                           from_latch_to_shifter_op1_9_port, a(8) => 
                           from_latch_to_shifter_op1_8_port, a(7) => 
                           from_latch_to_shifter_op1_7_port, a(6) => 
                           from_latch_to_shifter_op1_6_port, a(5) => 
                           from_latch_to_shifter_op1_5_port, a(4) => 
                           from_latch_to_shifter_op1_4_port, a(3) => 
                           from_latch_to_shifter_op1_3_port, a(2) => 
                           from_latch_to_shifter_op1_2_port, a(1) => 
                           from_latch_to_shifter_op1_1_port, a(0) => 
                           from_latch_to_shifter_op1_0_port, b(31) => 
                           from_latch_to_shifter_op2_31_port, b(30) => 
                           from_latch_to_shifter_op2_30_port, b(29) => 
                           from_latch_to_shifter_op2_29_port, b(28) => 
                           from_latch_to_shifter_op2_28_port, b(27) => 
                           from_latch_to_shifter_op2_27_port, b(26) => 
                           from_latch_to_shifter_op2_26_port, b(25) => 
                           from_latch_to_shifter_op2_25_port, b(24) => 
                           from_latch_to_shifter_op2_24_port, b(23) => 
                           from_latch_to_shifter_op2_23_port, b(22) => 
                           from_latch_to_shifter_op2_22_port, b(21) => 
                           from_latch_to_shifter_op2_21_port, b(20) => 
                           from_latch_to_shifter_op2_20_port, b(19) => 
                           from_latch_to_shifter_op2_19_port, b(18) => 
                           from_latch_to_shifter_op2_18_port, b(17) => 
                           from_latch_to_shifter_op2_17_port, b(16) => 
                           from_latch_to_shifter_op2_16_port, b(15) => 
                           from_latch_to_shifter_op2_15_port, b(14) => 
                           from_latch_to_shifter_op2_14_port, b(13) => 
                           from_latch_to_shifter_op2_13_port, b(12) => 
                           from_latch_to_shifter_op2_12_port, b(11) => 
                           from_latch_to_shifter_op2_11_port, b(10) => 
                           from_latch_to_shifter_op2_10_port, b(9) => 
                           from_latch_to_shifter_op2_9_port, b(8) => 
                           from_latch_to_shifter_op2_8_port, b(7) => 
                           from_latch_to_shifter_op2_7_port, b(6) => 
                           from_latch_to_shifter_op2_6_port, b(5) => 
                           from_latch_to_shifter_op2_5_port, b(4) => 
                           from_latch_to_shifter_op2_4_port, b(3) => 
                           from_latch_to_shifter_op2_3_port, b(2) => 
                           from_latch_to_shifter_op2_2_port, b(1) => 
                           from_latch_to_shifter_op2_1_port, b(0) => 
                           from_latch_to_shifter_op2_0_port, o(31) => 
                           from_shifter_to_mux_31_port, o(30) => 
                           from_shifter_to_mux_30_port, o(29) => 
                           from_shifter_to_mux_29_port, o(28) => 
                           from_shifter_to_mux_28_port, o(27) => 
                           from_shifter_to_mux_27_port, o(26) => 
                           from_shifter_to_mux_26_port, o(25) => 
                           from_shifter_to_mux_25_port, o(24) => 
                           from_shifter_to_mux_24_port, o(23) => 
                           from_shifter_to_mux_23_port, o(22) => 
                           from_shifter_to_mux_22_port, o(21) => 
                           from_shifter_to_mux_21_port, o(20) => 
                           from_shifter_to_mux_20_port, o(19) => 
                           from_shifter_to_mux_19_port, o(18) => 
                           from_shifter_to_mux_18_port, o(17) => 
                           from_shifter_to_mux_17_port, o(16) => 
                           from_shifter_to_mux_16_port, o(15) => 
                           from_shifter_to_mux_15_port, o(14) => 
                           from_shifter_to_mux_14_port, o(13) => 
                           from_shifter_to_mux_13_port, o(12) => 
                           from_shifter_to_mux_12_port, o(11) => 
                           from_shifter_to_mux_11_port, o(10) => 
                           from_shifter_to_mux_10_port, o(9) => 
                           from_shifter_to_mux_9_port, o(8) => 
                           from_shifter_to_mux_8_port, o(7) => 
                           from_shifter_to_mux_7_port, o(6) => 
                           from_shifter_to_mux_6_port, o(5) => 
                           from_shifter_to_mux_5_port, o(4) => 
                           from_shifter_to_mux_4_port, o(3) => 
                           from_shifter_to_mux_3_port, o(2) => 
                           from_shifter_to_mux_2_port, o(1) => 
                           from_shifter_to_mux_1_port, o(0) => 
                           from_shifter_to_mux_0_port);
   BM : booths_mul_N_bit16 port map( multiplier(15) => 
                           from_latch_to_mul_op2_15_port, multiplier(14) => 
                           from_latch_to_mul_op2_14_port, multiplier(13) => 
                           from_latch_to_mul_op2_13_port, multiplier(12) => 
                           from_latch_to_mul_op2_12_port, multiplier(11) => 
                           from_latch_to_mul_op2_11_port, multiplier(10) => 
                           from_latch_to_mul_op2_10_port, multiplier(9) => 
                           from_latch_to_mul_op2_9_port, multiplier(8) => 
                           from_latch_to_mul_op2_8_port, multiplier(7) => 
                           from_latch_to_mul_op2_7_port, multiplier(6) => 
                           from_latch_to_mul_op2_6_port, multiplier(5) => 
                           from_latch_to_mul_op2_5_port, multiplier(4) => 
                           from_latch_to_mul_op2_4_port, multiplier(3) => 
                           from_latch_to_mul_op2_3_port, multiplier(2) => 
                           from_latch_to_mul_op2_2_port, multiplier(1) => 
                           from_latch_to_mul_op2_1_port, multiplier(0) => 
                           from_latch_to_mul_op2_0_port, multiplicand(15) => 
                           from_latch_to_mul_op1_15_port, multiplicand(14) => 
                           from_latch_to_mul_op1_14_port, multiplicand(13) => 
                           from_latch_to_mul_op1_13_port, multiplicand(12) => 
                           from_latch_to_mul_op1_12_port, multiplicand(11) => 
                           from_latch_to_mul_op1_11_port, multiplicand(10) => 
                           from_latch_to_mul_op1_10_port, multiplicand(9) => 
                           from_latch_to_mul_op1_9_port, multiplicand(8) => 
                           from_latch_to_mul_op1_8_port, multiplicand(7) => 
                           from_latch_to_mul_op1_7_port, multiplicand(6) => 
                           from_latch_to_mul_op1_6_port, multiplicand(5) => 
                           from_latch_to_mul_op1_5_port, multiplicand(4) => 
                           from_latch_to_mul_op1_4_port, multiplicand(3) => 
                           from_latch_to_mul_op1_3_port, multiplicand(2) => 
                           from_latch_to_mul_op1_2_port, multiplicand(1) => 
                           from_latch_to_mul_op1_1_port, multiplicand(0) => 
                           from_latch_to_mul_op1_0_port, product(31) => 
                           from_mul_to_mux_31_port, product(30) => 
                           from_mul_to_mux_30_port, product(29) => 
                           from_mul_to_mux_29_port, product(28) => 
                           from_mul_to_mux_28_port, product(27) => 
                           from_mul_to_mux_27_port, product(26) => 
                           from_mul_to_mux_26_port, product(25) => 
                           from_mul_to_mux_25_port, product(24) => 
                           from_mul_to_mux_24_port, product(23) => 
                           from_mul_to_mux_23_port, product(22) => 
                           from_mul_to_mux_22_port, product(21) => 
                           from_mul_to_mux_21_port, product(20) => 
                           from_mul_to_mux_20_port, product(19) => 
                           from_mul_to_mux_19_port, product(18) => 
                           from_mul_to_mux_18_port, product(17) => 
                           from_mul_to_mux_17_port, product(16) => 
                           from_mul_to_mux_16_port, product(15) => 
                           from_mul_to_mux_15_port, product(14) => 
                           from_mul_to_mux_14_port, product(13) => 
                           from_mul_to_mux_13_port, product(12) => 
                           from_mul_to_mux_12_port, product(11) => 
                           from_mul_to_mux_11_port, product(10) => 
                           from_mul_to_mux_10_port, product(9) => 
                           from_mul_to_mux_9_port, product(8) => 
                           from_mul_to_mux_8_port, product(7) => 
                           from_mul_to_mux_7_port, product(6) => 
                           from_mul_to_mux_6_port, product(5) => 
                           from_mul_to_mux_5_port, product(4) => 
                           from_mul_to_mux_4_port, product(3) => 
                           from_mul_to_mux_3_port, product(2) => 
                           from_mul_to_mux_2_port, product(1) => 
                           from_mul_to_mux_1_port, product(0) => 
                           from_mul_to_mux_0_port);
   M4 : mux5x1 port map( a(31) => from_adder_to_mux_31_port, a(30) => 
                           from_adder_to_mux_30_port, a(29) => 
                           from_adder_to_mux_29_port, a(28) => 
                           from_adder_to_mux_28_port, a(27) => 
                           from_adder_to_mux_27_port, a(26) => 
                           from_adder_to_mux_26_port, a(25) => 
                           from_adder_to_mux_25_port, a(24) => 
                           from_adder_to_mux_24_port, a(23) => 
                           from_adder_to_mux_23_port, a(22) => 
                           from_adder_to_mux_22_port, a(21) => 
                           from_adder_to_mux_21_port, a(20) => 
                           from_adder_to_mux_20_port, a(19) => 
                           from_adder_to_mux_19_port, a(18) => 
                           from_adder_to_mux_18_port, a(17) => 
                           from_adder_to_mux_17_port, a(16) => 
                           from_adder_to_mux_16_port, a(15) => 
                           from_adder_to_mux_15_port, a(14) => 
                           from_adder_to_mux_14_port, a(13) => 
                           from_adder_to_mux_13_port, a(12) => 
                           from_adder_to_mux_12_port, a(11) => 
                           from_adder_to_mux_11_port, a(10) => 
                           from_adder_to_mux_10_port, a(9) => 
                           from_adder_to_mux_9_port, a(8) => 
                           from_adder_to_mux_8_port, a(7) => 
                           from_adder_to_mux_7_port, a(6) => 
                           from_adder_to_mux_6_port, a(5) => 
                           from_adder_to_mux_5_port, a(4) => 
                           from_adder_to_mux_4_port, a(3) => 
                           from_adder_to_mux_3_port, a(2) => 
                           from_adder_to_mux_2_port, a(1) => 
                           from_adder_to_mux_1_port, a(0) => 
                           from_adder_to_mux_0_port, b(31) => 
                           from_logict2_to_mux_31_port, b(30) => 
                           from_logict2_to_mux_30_port, b(29) => 
                           from_logict2_to_mux_29_port, b(28) => 
                           from_logict2_to_mux_28_port, b(27) => 
                           from_logict2_to_mux_27_port, b(26) => 
                           from_logict2_to_mux_26_port, b(25) => 
                           from_logict2_to_mux_25_port, b(24) => 
                           from_logict2_to_mux_24_port, b(23) => 
                           from_logict2_to_mux_23_port, b(22) => 
                           from_logict2_to_mux_22_port, b(21) => 
                           from_logict2_to_mux_21_port, b(20) => 
                           from_logict2_to_mux_20_port, b(19) => 
                           from_logict2_to_mux_19_port, b(18) => 
                           from_logict2_to_mux_18_port, b(17) => 
                           from_logict2_to_mux_17_port, b(16) => 
                           from_logict2_to_mux_16_port, b(15) => 
                           from_logict2_to_mux_15_port, b(14) => 
                           from_logict2_to_mux_14_port, b(13) => 
                           from_logict2_to_mux_13_port, b(12) => 
                           from_logict2_to_mux_12_port, b(11) => 
                           from_logict2_to_mux_11_port, b(10) => 
                           from_logict2_to_mux_10_port, b(9) => 
                           from_logict2_to_mux_9_port, b(8) => 
                           from_logict2_to_mux_8_port, b(7) => 
                           from_logict2_to_mux_7_port, b(6) => 
                           from_logict2_to_mux_6_port, b(5) => 
                           from_logict2_to_mux_5_port, b(4) => 
                           from_logict2_to_mux_4_port, b(3) => 
                           from_logict2_to_mux_3_port, b(2) => 
                           from_logict2_to_mux_2_port, b(1) => 
                           from_logict2_to_mux_1_port, b(0) => 
                           from_logict2_to_mux_0_port, c(31) => 
                           from_mul_to_mux_31_port, c(30) => 
                           from_mul_to_mux_30_port, c(29) => 
                           from_mul_to_mux_29_port, c(28) => 
                           from_mul_to_mux_28_port, c(27) => 
                           from_mul_to_mux_27_port, c(26) => 
                           from_mul_to_mux_26_port, c(25) => 
                           from_mul_to_mux_25_port, c(24) => 
                           from_mul_to_mux_24_port, c(23) => 
                           from_mul_to_mux_23_port, c(22) => 
                           from_mul_to_mux_22_port, c(21) => 
                           from_mul_to_mux_21_port, c(20) => 
                           from_mul_to_mux_20_port, c(19) => 
                           from_mul_to_mux_19_port, c(18) => 
                           from_mul_to_mux_18_port, c(17) => 
                           from_mul_to_mux_17_port, c(16) => 
                           from_mul_to_mux_16_port, c(15) => 
                           from_mul_to_mux_15_port, c(14) => 
                           from_mul_to_mux_14_port, c(13) => 
                           from_mul_to_mux_13_port, c(12) => 
                           from_mul_to_mux_12_port, c(11) => 
                           from_mul_to_mux_11_port, c(10) => 
                           from_mul_to_mux_10_port, c(9) => 
                           from_mul_to_mux_9_port, c(8) => 
                           from_mul_to_mux_8_port, c(7) => 
                           from_mul_to_mux_7_port, c(6) => 
                           from_mul_to_mux_6_port, c(5) => 
                           from_mul_to_mux_5_port, c(4) => 
                           from_mul_to_mux_4_port, c(3) => 
                           from_mul_to_mux_3_port, c(2) => 
                           from_mul_to_mux_2_port, c(1) => 
                           from_mul_to_mux_1_port, c(0) => 
                           from_mul_to_mux_0_port, d(31) => 
                           from_shifter_to_mux_31_port, d(30) => 
                           from_shifter_to_mux_30_port, d(29) => 
                           from_shifter_to_mux_29_port, d(28) => 
                           from_shifter_to_mux_28_port, d(27) => 
                           from_shifter_to_mux_27_port, d(26) => 
                           from_shifter_to_mux_26_port, d(25) => 
                           from_shifter_to_mux_25_port, d(24) => 
                           from_shifter_to_mux_24_port, d(23) => 
                           from_shifter_to_mux_23_port, d(22) => 
                           from_shifter_to_mux_22_port, d(21) => 
                           from_shifter_to_mux_21_port, d(20) => 
                           from_shifter_to_mux_20_port, d(19) => 
                           from_shifter_to_mux_19_port, d(18) => 
                           from_shifter_to_mux_18_port, d(17) => 
                           from_shifter_to_mux_17_port, d(16) => 
                           from_shifter_to_mux_16_port, d(15) => 
                           from_shifter_to_mux_15_port, d(14) => 
                           from_shifter_to_mux_14_port, d(13) => 
                           from_shifter_to_mux_13_port, d(12) => 
                           from_shifter_to_mux_12_port, d(11) => 
                           from_shifter_to_mux_11_port, d(10) => 
                           from_shifter_to_mux_10_port, d(9) => 
                           from_shifter_to_mux_9_port, d(8) => 
                           from_shifter_to_mux_8_port, d(7) => 
                           from_shifter_to_mux_7_port, d(6) => 
                           from_shifter_to_mux_6_port, d(5) => 
                           from_shifter_to_mux_5_port, d(4) => 
                           from_shifter_to_mux_4_port, d(3) => 
                           from_shifter_to_mux_3_port, d(2) => 
                           from_shifter_to_mux_2_port, d(1) => 
                           from_shifter_to_mux_1_port, d(0) => 
                           from_shifter_to_mux_0_port, e(31) => 
                           from_comparator_to_mux_31_port, e(30) => 
                           from_comparator_to_mux_30_port, e(29) => 
                           from_comparator_to_mux_29_port, e(28) => 
                           from_comparator_to_mux_28_port, e(27) => 
                           from_comparator_to_mux_27_port, e(26) => 
                           from_comparator_to_mux_26_port, e(25) => 
                           from_comparator_to_mux_25_port, e(24) => 
                           from_comparator_to_mux_24_port, e(23) => 
                           from_comparator_to_mux_23_port, e(22) => 
                           from_comparator_to_mux_22_port, e(21) => 
                           from_comparator_to_mux_21_port, e(20) => 
                           from_comparator_to_mux_20_port, e(19) => 
                           from_comparator_to_mux_19_port, e(18) => 
                           from_comparator_to_mux_18_port, e(17) => 
                           from_comparator_to_mux_17_port, e(16) => 
                           from_comparator_to_mux_16_port, e(15) => 
                           from_comparator_to_mux_15_port, e(14) => 
                           from_comparator_to_mux_14_port, e(13) => 
                           from_comparator_to_mux_13_port, e(12) => 
                           from_comparator_to_mux_12_port, e(11) => 
                           from_comparator_to_mux_11_port, e(10) => 
                           from_comparator_to_mux_10_port, e(9) => 
                           from_comparator_to_mux_9_port, e(8) => 
                           from_comparator_to_mux_8_port, e(7) => 
                           from_comparator_to_mux_7_port, e(6) => 
                           from_comparator_to_mux_6_port, e(5) => 
                           from_comparator_to_mux_5_port, e(4) => 
                           from_comparator_to_mux_4_port, e(3) => 
                           from_comparator_to_mux_3_port, e(2) => 
                           from_comparator_to_mux_2_port, e(1) => 
                           from_comparator_to_mux_1_port, e(0) => jump_port, 
                           enable => enable_mux_4_1, sel(2) => 
                           sel_signal_5_1_2_port, sel(1) => 
                           sel_signal_5_1_1_port, sel(0) => 
                           sel_signal_5_1_0_port, out_res(31) => 
                           from_mux_4_1_to_mux_2_1_31_port, out_res(30) => 
                           from_mux_4_1_to_mux_2_1_30_port, out_res(29) => 
                           from_mux_4_1_to_mux_2_1_29_port, out_res(28) => 
                           from_mux_4_1_to_mux_2_1_28_port, out_res(27) => 
                           from_mux_4_1_to_mux_2_1_27_port, out_res(26) => 
                           from_mux_4_1_to_mux_2_1_26_port, out_res(25) => 
                           from_mux_4_1_to_mux_2_1_25_port, out_res(24) => 
                           from_mux_4_1_to_mux_2_1_24_port, out_res(23) => 
                           from_mux_4_1_to_mux_2_1_23_port, out_res(22) => 
                           from_mux_4_1_to_mux_2_1_22_port, out_res(21) => 
                           from_mux_4_1_to_mux_2_1_21_port, out_res(20) => 
                           from_mux_4_1_to_mux_2_1_20_port, out_res(19) => 
                           from_mux_4_1_to_mux_2_1_19_port, out_res(18) => 
                           from_mux_4_1_to_mux_2_1_18_port, out_res(17) => 
                           from_mux_4_1_to_mux_2_1_17_port, out_res(16) => 
                           from_mux_4_1_to_mux_2_1_16_port, out_res(15) => 
                           from_mux_4_1_to_mux_2_1_15_port, out_res(14) => 
                           from_mux_4_1_to_mux_2_1_14_port, out_res(13) => 
                           from_mux_4_1_to_mux_2_1_13_port, out_res(12) => 
                           from_mux_4_1_to_mux_2_1_12_port, out_res(11) => 
                           from_mux_4_1_to_mux_2_1_11_port, out_res(10) => 
                           from_mux_4_1_to_mux_2_1_10_port, out_res(9) => 
                           from_mux_4_1_to_mux_2_1_9_port, out_res(8) => 
                           from_mux_4_1_to_mux_2_1_8_port, out_res(7) => 
                           from_mux_4_1_to_mux_2_1_7_port, out_res(6) => 
                           from_mux_4_1_to_mux_2_1_6_port, out_res(5) => 
                           from_mux_4_1_to_mux_2_1_5_port, out_res(4) => 
                           from_mux_4_1_to_mux_2_1_4_port, out_res(3) => 
                           from_mux_4_1_to_mux_2_1_3_port, out_res(2) => 
                           from_mux_4_1_to_mux_2_1_2_port, out_res(1) => 
                           from_mux_4_1_to_mux_2_1_1_port, out_res(0) => 
                           from_mux_4_1_to_mux_2_1_0_port);
   T2 : logicUnitT2_data_size32 port map( operand_a(31) => 
                           from_latch_to_logict2_op1_31_port, operand_a(30) => 
                           from_latch_to_logict2_op1_30_port, operand_a(29) => 
                           from_latch_to_logict2_op1_29_port, operand_a(28) => 
                           from_latch_to_logict2_op1_28_port, operand_a(27) => 
                           from_latch_to_logict2_op1_27_port, operand_a(26) => 
                           from_latch_to_logict2_op1_26_port, operand_a(25) => 
                           from_latch_to_logict2_op1_25_port, operand_a(24) => 
                           from_latch_to_logict2_op1_24_port, operand_a(23) => 
                           from_latch_to_logict2_op1_23_port, operand_a(22) => 
                           from_latch_to_logict2_op1_22_port, operand_a(21) => 
                           from_latch_to_logict2_op1_21_port, operand_a(20) => 
                           from_latch_to_logict2_op1_20_port, operand_a(19) => 
                           from_latch_to_logict2_op1_19_port, operand_a(18) => 
                           from_latch_to_logict2_op1_18_port, operand_a(17) => 
                           from_latch_to_logict2_op1_17_port, operand_a(16) => 
                           from_latch_to_logict2_op1_16_port, operand_a(15) => 
                           from_latch_to_logict2_op1_15_port, operand_a(14) => 
                           from_latch_to_logict2_op1_14_port, operand_a(13) => 
                           from_latch_to_logict2_op1_13_port, operand_a(12) => 
                           from_latch_to_logict2_op1_12_port, operand_a(11) => 
                           from_latch_to_logict2_op1_11_port, operand_a(10) => 
                           from_latch_to_logict2_op1_10_port, operand_a(9) => 
                           from_latch_to_logict2_op1_9_port, operand_a(8) => 
                           from_latch_to_logict2_op1_8_port, operand_a(7) => 
                           from_latch_to_logict2_op1_7_port, operand_a(6) => 
                           from_latch_to_logict2_op1_6_port, operand_a(5) => 
                           from_latch_to_logict2_op1_5_port, operand_a(4) => 
                           from_latch_to_logict2_op1_4_port, operand_a(3) => 
                           from_latch_to_logict2_op1_3_port, operand_a(2) => 
                           from_latch_to_logict2_op1_2_port, operand_a(1) => 
                           from_latch_to_logict2_op1_1_port, operand_a(0) => 
                           from_latch_to_logict2_op1_0_port, operand_b(31) => 
                           from_latch_to_logict2_op2_31_port, operand_b(30) => 
                           from_latch_to_logict2_op2_30_port, operand_b(29) => 
                           from_latch_to_logict2_op2_29_port, operand_b(28) => 
                           from_latch_to_logict2_op2_28_port, operand_b(27) => 
                           from_latch_to_logict2_op2_27_port, operand_b(26) => 
                           from_latch_to_logict2_op2_26_port, operand_b(25) => 
                           from_latch_to_logict2_op2_25_port, operand_b(24) => 
                           from_latch_to_logict2_op2_24_port, operand_b(23) => 
                           from_latch_to_logict2_op2_23_port, operand_b(22) => 
                           from_latch_to_logict2_op2_22_port, operand_b(21) => 
                           from_latch_to_logict2_op2_21_port, operand_b(20) => 
                           from_latch_to_logict2_op2_20_port, operand_b(19) => 
                           from_latch_to_logict2_op2_19_port, operand_b(18) => 
                           from_latch_to_logict2_op2_18_port, operand_b(17) => 
                           from_latch_to_logict2_op2_17_port, operand_b(16) => 
                           from_latch_to_logict2_op2_16_port, operand_b(15) => 
                           from_latch_to_logict2_op2_15_port, operand_b(14) => 
                           from_latch_to_logict2_op2_14_port, operand_b(13) => 
                           from_latch_to_logict2_op2_13_port, operand_b(12) => 
                           from_latch_to_logict2_op2_12_port, operand_b(11) => 
                           from_latch_to_logict2_op2_11_port, operand_b(10) => 
                           from_latch_to_logict2_op2_10_port, operand_b(9) => 
                           from_latch_to_logict2_op2_9_port, operand_b(8) => 
                           from_latch_to_logict2_op2_8_port, operand_b(7) => 
                           from_latch_to_logict2_op2_7_port, operand_b(6) => 
                           from_latch_to_logict2_op2_6_port, operand_b(5) => 
                           from_latch_to_logict2_op2_5_port, operand_b(4) => 
                           from_latch_to_logict2_op2_4_port, operand_b(3) => 
                           from_latch_to_logict2_op2_3_port, operand_b(2) => 
                           from_latch_to_logict2_op2_2_port, operand_b(1) => 
                           from_latch_to_logict2_op2_1_port, operand_b(0) => 
                           from_latch_to_logict2_op2_0_port, type_op(3) => 
                           signal_cmd_t2_3_port, type_op(2) => 
                           signal_cmd_t2_2_port, type_op(1) => 
                           signal_cmd_t2_1_port, type_op(0) => 
                           signal_cmd_t2_0_port, result(31) => 
                           from_logict2_to_mux_31_port, result(30) => 
                           from_logict2_to_mux_30_port, result(29) => 
                           from_logict2_to_mux_29_port, result(28) => 
                           from_logict2_to_mux_28_port, result(27) => 
                           from_logict2_to_mux_27_port, result(26) => 
                           from_logict2_to_mux_26_port, result(25) => 
                           from_logict2_to_mux_25_port, result(24) => 
                           from_logict2_to_mux_24_port, result(23) => 
                           from_logict2_to_mux_23_port, result(22) => 
                           from_logict2_to_mux_22_port, result(21) => 
                           from_logict2_to_mux_21_port, result(20) => 
                           from_logict2_to_mux_20_port, result(19) => 
                           from_logict2_to_mux_19_port, result(18) => 
                           from_logict2_to_mux_18_port, result(17) => 
                           from_logict2_to_mux_17_port, result(16) => 
                           from_logict2_to_mux_16_port, result(15) => 
                           from_logict2_to_mux_15_port, result(14) => 
                           from_logict2_to_mux_14_port, result(13) => 
                           from_logict2_to_mux_13_port, result(12) => 
                           from_logict2_to_mux_12_port, result(11) => 
                           from_logict2_to_mux_11_port, result(10) => 
                           from_logict2_to_mux_10_port, result(9) => 
                           from_logict2_to_mux_9_port, result(8) => 
                           from_logict2_to_mux_8_port, result(7) => 
                           from_logict2_to_mux_7_port, result(6) => 
                           from_logict2_to_mux_6_port, result(5) => 
                           from_logict2_to_mux_5_port, result(4) => 
                           from_logict2_to_mux_4_port, result(3) => 
                           from_logict2_to_mux_3_port, result(2) => 
                           from_logict2_to_mux_2_port, result(1) => 
                           from_logict2_to_mux_1_port, result(0) => 
                           from_logict2_to_mux_0_port);
   PL0 : positive_latch_on_000_0 port map( d(31) => 
                           from_mux_2_1_to_latch_high_31_port, d(30) => 
                           from_mux_2_1_to_latch_high_30_port, d(29) => 
                           from_mux_2_1_to_latch_high_29_port, d(28) => 
                           from_mux_2_1_to_latch_high_28_port, d(27) => 
                           from_mux_2_1_to_latch_high_27_port, d(26) => 
                           from_mux_2_1_to_latch_high_26_port, d(25) => 
                           from_mux_2_1_to_latch_high_25_port, d(24) => 
                           from_mux_2_1_to_latch_high_24_port, d(23) => 
                           from_mux_2_1_to_latch_high_23_port, d(22) => 
                           from_mux_2_1_to_latch_high_22_port, d(21) => 
                           from_mux_2_1_to_latch_high_21_port, d(20) => 
                           from_mux_2_1_to_latch_high_20_port, d(19) => 
                           from_mux_2_1_to_latch_high_19_port, d(18) => 
                           from_mux_2_1_to_latch_high_18_port, d(17) => 
                           from_mux_2_1_to_latch_high_17_port, d(16) => 
                           from_mux_2_1_to_latch_high_16_port, d(15) => 
                           from_mux_2_1_to_latch_high_15_port, d(14) => 
                           from_mux_2_1_to_latch_high_14_port, d(13) => 
                           from_mux_2_1_to_latch_high_13_port, d(12) => 
                           from_mux_2_1_to_latch_high_12_port, d(11) => 
                           from_mux_2_1_to_latch_high_11_port, d(10) => 
                           from_mux_2_1_to_latch_high_10_port, d(9) => 
                           from_mux_2_1_to_latch_high_9_port, d(8) => 
                           from_mux_2_1_to_latch_high_8_port, d(7) => 
                           from_mux_2_1_to_latch_high_7_port, d(6) => 
                           from_mux_2_1_to_latch_high_6_port, d(5) => 
                           from_mux_2_1_to_latch_high_5_port, d(4) => 
                           from_mux_2_1_to_latch_high_4_port, d(3) => 
                           from_mux_2_1_to_latch_high_3_port, d(2) => 
                           from_mux_2_1_to_latch_high_2_port, d(1) => 
                           from_mux_2_1_to_latch_high_1_port, d(0) => 
                           from_mux_2_1_to_latch_high_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_adder_op1_31_port, q(30) => 
                           from_latch_to_adder_op1_30_port, q(29) => 
                           from_latch_to_adder_op1_29_port, q(28) => 
                           from_latch_to_adder_op1_28_port, q(27) => 
                           from_latch_to_adder_op1_27_port, q(26) => 
                           from_latch_to_adder_op1_26_port, q(25) => 
                           from_latch_to_adder_op1_25_port, q(24) => 
                           from_latch_to_adder_op1_24_port, q(23) => 
                           from_latch_to_adder_op1_23_port, q(22) => 
                           from_latch_to_adder_op1_22_port, q(21) => 
                           from_latch_to_adder_op1_21_port, q(20) => 
                           from_latch_to_adder_op1_20_port, q(19) => 
                           from_latch_to_adder_op1_19_port, q(18) => 
                           from_latch_to_adder_op1_18_port, q(17) => 
                           from_latch_to_adder_op1_17_port, q(16) => 
                           from_latch_to_adder_op1_16_port, q(15) => 
                           from_latch_to_adder_op1_15_port, q(14) => 
                           from_latch_to_adder_op1_14_port, q(13) => 
                           from_latch_to_adder_op1_13_port, q(12) => 
                           from_latch_to_adder_op1_12_port, q(11) => 
                           from_latch_to_adder_op1_11_port, q(10) => 
                           from_latch_to_adder_op1_10_port, q(9) => 
                           from_latch_to_adder_op1_9_port, q(8) => 
                           from_latch_to_adder_op1_8_port, q(7) => 
                           from_latch_to_adder_op1_7_port, q(6) => 
                           from_latch_to_adder_op1_6_port, q(5) => 
                           from_latch_to_adder_op1_5_port, q(4) => 
                           from_latch_to_adder_op1_4_port, q(3) => 
                           from_latch_to_adder_op1_3_port, q(2) => 
                           from_latch_to_adder_op1_2_port, q(1) => 
                           from_latch_to_adder_op1_1_port, q(0) => 
                           from_latch_to_adder_op1_0_port);
   PL1 : positive_latch_on_000_1 port map( d(31) => 
                           from_mux_2_1_to_latch_low_31_port, d(30) => 
                           from_mux_2_1_to_latch_low_30_port, d(29) => 
                           from_mux_2_1_to_latch_low_29_port, d(28) => 
                           from_mux_2_1_to_latch_low_28_port, d(27) => 
                           from_mux_2_1_to_latch_low_27_port, d(26) => 
                           from_mux_2_1_to_latch_low_26_port, d(25) => 
                           from_mux_2_1_to_latch_low_25_port, d(24) => 
                           from_mux_2_1_to_latch_low_24_port, d(23) => 
                           from_mux_2_1_to_latch_low_23_port, d(22) => 
                           from_mux_2_1_to_latch_low_22_port, d(21) => 
                           from_mux_2_1_to_latch_low_21_port, d(20) => 
                           from_mux_2_1_to_latch_low_20_port, d(19) => 
                           from_mux_2_1_to_latch_low_19_port, d(18) => 
                           from_mux_2_1_to_latch_low_18_port, d(17) => 
                           from_mux_2_1_to_latch_low_17_port, d(16) => 
                           from_mux_2_1_to_latch_low_16_port, d(15) => 
                           from_mux_2_1_to_latch_low_15_port, d(14) => 
                           from_mux_2_1_to_latch_low_14_port, d(13) => 
                           from_mux_2_1_to_latch_low_13_port, d(12) => 
                           from_mux_2_1_to_latch_low_12_port, d(11) => 
                           from_mux_2_1_to_latch_low_11_port, d(10) => 
                           from_mux_2_1_to_latch_low_10_port, d(9) => 
                           from_mux_2_1_to_latch_low_9_port, d(8) => 
                           from_mux_2_1_to_latch_low_8_port, d(7) => 
                           from_mux_2_1_to_latch_low_7_port, d(6) => 
                           from_mux_2_1_to_latch_low_6_port, d(5) => 
                           from_mux_2_1_to_latch_low_5_port, d(4) => 
                           from_mux_2_1_to_latch_low_4_port, d(3) => 
                           from_mux_2_1_to_latch_low_3_port, d(2) => 
                           from_mux_2_1_to_latch_low_2_port, d(1) => 
                           from_mux_2_1_to_latch_low_1_port, d(0) => 
                           from_mux_2_1_to_latch_low_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_mux_sub_or_add_31_port, q(30) => 
                           from_latch_to_mux_sub_or_add_30_port, q(29) => 
                           from_latch_to_mux_sub_or_add_29_port, q(28) => 
                           from_latch_to_mux_sub_or_add_28_port, q(27) => 
                           from_latch_to_mux_sub_or_add_27_port, q(26) => 
                           from_latch_to_mux_sub_or_add_26_port, q(25) => 
                           from_latch_to_mux_sub_or_add_25_port, q(24) => 
                           from_latch_to_mux_sub_or_add_24_port, q(23) => 
                           from_latch_to_mux_sub_or_add_23_port, q(22) => 
                           from_latch_to_mux_sub_or_add_22_port, q(21) => 
                           from_latch_to_mux_sub_or_add_21_port, q(20) => 
                           from_latch_to_mux_sub_or_add_20_port, q(19) => 
                           from_latch_to_mux_sub_or_add_19_port, q(18) => 
                           from_latch_to_mux_sub_or_add_18_port, q(17) => 
                           from_latch_to_mux_sub_or_add_17_port, q(16) => 
                           from_latch_to_mux_sub_or_add_16_port, q(15) => 
                           from_latch_to_mux_sub_or_add_15_port, q(14) => 
                           from_latch_to_mux_sub_or_add_14_port, q(13) => 
                           from_latch_to_mux_sub_or_add_13_port, q(12) => 
                           from_latch_to_mux_sub_or_add_12_port, q(11) => 
                           from_latch_to_mux_sub_or_add_11_port, q(10) => 
                           from_latch_to_mux_sub_or_add_10_port, q(9) => 
                           from_latch_to_mux_sub_or_add_9_port, q(8) => 
                           from_latch_to_mux_sub_or_add_8_port, q(7) => 
                           from_latch_to_mux_sub_or_add_7_port, q(6) => 
                           from_latch_to_mux_sub_or_add_6_port, q(5) => 
                           from_latch_to_mux_sub_or_add_5_port, q(4) => 
                           from_latch_to_mux_sub_or_add_4_port, q(3) => 
                           from_latch_to_mux_sub_or_add_3_port, q(2) => 
                           from_latch_to_mux_sub_or_add_2_port, q(1) => 
                           from_latch_to_mux_sub_or_add_1_port, q(0) => 
                           from_latch_to_mux_sub_or_add_0_port);
   PL2 : positive_latch_on_001_0 port map( d(31) => 
                           from_mux_2_1_to_latch_high_31_port, d(30) => 
                           from_mux_2_1_to_latch_high_30_port, d(29) => 
                           from_mux_2_1_to_latch_high_29_port, d(28) => 
                           from_mux_2_1_to_latch_high_28_port, d(27) => 
                           from_mux_2_1_to_latch_high_27_port, d(26) => 
                           from_mux_2_1_to_latch_high_26_port, d(25) => 
                           from_mux_2_1_to_latch_high_25_port, d(24) => 
                           from_mux_2_1_to_latch_high_24_port, d(23) => 
                           from_mux_2_1_to_latch_high_23_port, d(22) => 
                           from_mux_2_1_to_latch_high_22_port, d(21) => 
                           from_mux_2_1_to_latch_high_21_port, d(20) => 
                           from_mux_2_1_to_latch_high_20_port, d(19) => 
                           from_mux_2_1_to_latch_high_19_port, d(18) => 
                           from_mux_2_1_to_latch_high_18_port, d(17) => 
                           from_mux_2_1_to_latch_high_17_port, d(16) => 
                           from_mux_2_1_to_latch_high_16_port, d(15) => 
                           from_mux_2_1_to_latch_high_15_port, d(14) => 
                           from_mux_2_1_to_latch_high_14_port, d(13) => 
                           from_mux_2_1_to_latch_high_13_port, d(12) => 
                           from_mux_2_1_to_latch_high_12_port, d(11) => 
                           from_mux_2_1_to_latch_high_11_port, d(10) => 
                           from_mux_2_1_to_latch_high_10_port, d(9) => 
                           from_mux_2_1_to_latch_high_9_port, d(8) => 
                           from_mux_2_1_to_latch_high_8_port, d(7) => 
                           from_mux_2_1_to_latch_high_7_port, d(6) => 
                           from_mux_2_1_to_latch_high_6_port, d(5) => 
                           from_mux_2_1_to_latch_high_5_port, d(4) => 
                           from_mux_2_1_to_latch_high_4_port, d(3) => 
                           from_mux_2_1_to_latch_high_3_port, d(2) => 
                           from_mux_2_1_to_latch_high_2_port, d(1) => 
                           from_mux_2_1_to_latch_high_1_port, d(0) => 
                           from_mux_2_1_to_latch_high_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_logict2_op1_31_port, q(30) => 
                           from_latch_to_logict2_op1_30_port, q(29) => 
                           from_latch_to_logict2_op1_29_port, q(28) => 
                           from_latch_to_logict2_op1_28_port, q(27) => 
                           from_latch_to_logict2_op1_27_port, q(26) => 
                           from_latch_to_logict2_op1_26_port, q(25) => 
                           from_latch_to_logict2_op1_25_port, q(24) => 
                           from_latch_to_logict2_op1_24_port, q(23) => 
                           from_latch_to_logict2_op1_23_port, q(22) => 
                           from_latch_to_logict2_op1_22_port, q(21) => 
                           from_latch_to_logict2_op1_21_port, q(20) => 
                           from_latch_to_logict2_op1_20_port, q(19) => 
                           from_latch_to_logict2_op1_19_port, q(18) => 
                           from_latch_to_logict2_op1_18_port, q(17) => 
                           from_latch_to_logict2_op1_17_port, q(16) => 
                           from_latch_to_logict2_op1_16_port, q(15) => 
                           from_latch_to_logict2_op1_15_port, q(14) => 
                           from_latch_to_logict2_op1_14_port, q(13) => 
                           from_latch_to_logict2_op1_13_port, q(12) => 
                           from_latch_to_logict2_op1_12_port, q(11) => 
                           from_latch_to_logict2_op1_11_port, q(10) => 
                           from_latch_to_logict2_op1_10_port, q(9) => 
                           from_latch_to_logict2_op1_9_port, q(8) => 
                           from_latch_to_logict2_op1_8_port, q(7) => 
                           from_latch_to_logict2_op1_7_port, q(6) => 
                           from_latch_to_logict2_op1_6_port, q(5) => 
                           from_latch_to_logict2_op1_5_port, q(4) => 
                           from_latch_to_logict2_op1_4_port, q(3) => 
                           from_latch_to_logict2_op1_3_port, q(2) => 
                           from_latch_to_logict2_op1_2_port, q(1) => 
                           from_latch_to_logict2_op1_1_port, q(0) => 
                           from_latch_to_logict2_op1_0_port);
   PL3 : positive_latch_on_001_1 port map( d(31) => 
                           from_mux_2_1_to_latch_low_31_port, d(30) => 
                           from_mux_2_1_to_latch_low_30_port, d(29) => 
                           from_mux_2_1_to_latch_low_29_port, d(28) => 
                           from_mux_2_1_to_latch_low_28_port, d(27) => 
                           from_mux_2_1_to_latch_low_27_port, d(26) => 
                           from_mux_2_1_to_latch_low_26_port, d(25) => 
                           from_mux_2_1_to_latch_low_25_port, d(24) => 
                           from_mux_2_1_to_latch_low_24_port, d(23) => 
                           from_mux_2_1_to_latch_low_23_port, d(22) => 
                           from_mux_2_1_to_latch_low_22_port, d(21) => 
                           from_mux_2_1_to_latch_low_21_port, d(20) => 
                           from_mux_2_1_to_latch_low_20_port, d(19) => 
                           from_mux_2_1_to_latch_low_19_port, d(18) => 
                           from_mux_2_1_to_latch_low_18_port, d(17) => 
                           from_mux_2_1_to_latch_low_17_port, d(16) => 
                           from_mux_2_1_to_latch_low_16_port, d(15) => 
                           from_mux_2_1_to_latch_low_15_port, d(14) => 
                           from_mux_2_1_to_latch_low_14_port, d(13) => 
                           from_mux_2_1_to_latch_low_13_port, d(12) => 
                           from_mux_2_1_to_latch_low_12_port, d(11) => 
                           from_mux_2_1_to_latch_low_11_port, d(10) => 
                           from_mux_2_1_to_latch_low_10_port, d(9) => 
                           from_mux_2_1_to_latch_low_9_port, d(8) => 
                           from_mux_2_1_to_latch_low_8_port, d(7) => 
                           from_mux_2_1_to_latch_low_7_port, d(6) => 
                           from_mux_2_1_to_latch_low_6_port, d(5) => 
                           from_mux_2_1_to_latch_low_5_port, d(4) => 
                           from_mux_2_1_to_latch_low_4_port, d(3) => 
                           from_mux_2_1_to_latch_low_3_port, d(2) => 
                           from_mux_2_1_to_latch_low_2_port, d(1) => 
                           from_mux_2_1_to_latch_low_1_port, d(0) => 
                           from_mux_2_1_to_latch_low_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_logict2_op2_31_port, q(30) => 
                           from_latch_to_logict2_op2_30_port, q(29) => 
                           from_latch_to_logict2_op2_29_port, q(28) => 
                           from_latch_to_logict2_op2_28_port, q(27) => 
                           from_latch_to_logict2_op2_27_port, q(26) => 
                           from_latch_to_logict2_op2_26_port, q(25) => 
                           from_latch_to_logict2_op2_25_port, q(24) => 
                           from_latch_to_logict2_op2_24_port, q(23) => 
                           from_latch_to_logict2_op2_23_port, q(22) => 
                           from_latch_to_logict2_op2_22_port, q(21) => 
                           from_latch_to_logict2_op2_21_port, q(20) => 
                           from_latch_to_logict2_op2_20_port, q(19) => 
                           from_latch_to_logict2_op2_19_port, q(18) => 
                           from_latch_to_logict2_op2_18_port, q(17) => 
                           from_latch_to_logict2_op2_17_port, q(16) => 
                           from_latch_to_logict2_op2_16_port, q(15) => 
                           from_latch_to_logict2_op2_15_port, q(14) => 
                           from_latch_to_logict2_op2_14_port, q(13) => 
                           from_latch_to_logict2_op2_13_port, q(12) => 
                           from_latch_to_logict2_op2_12_port, q(11) => 
                           from_latch_to_logict2_op2_11_port, q(10) => 
                           from_latch_to_logict2_op2_10_port, q(9) => 
                           from_latch_to_logict2_op2_9_port, q(8) => 
                           from_latch_to_logict2_op2_8_port, q(7) => 
                           from_latch_to_logict2_op2_7_port, q(6) => 
                           from_latch_to_logict2_op2_6_port, q(5) => 
                           from_latch_to_logict2_op2_5_port, q(4) => 
                           from_latch_to_logict2_op2_4_port, q(3) => 
                           from_latch_to_logict2_op2_3_port, q(2) => 
                           from_latch_to_logict2_op2_2_port, q(1) => 
                           from_latch_to_logict2_op2_1_port, q(0) => 
                           from_latch_to_logict2_op2_0_port);
   PL4 : positive_latch_on_010_0 port map( d(31) => 
                           from_mux_2_1_to_latch_high_31_port, d(30) => 
                           from_mux_2_1_to_latch_high_30_port, d(29) => 
                           from_mux_2_1_to_latch_high_29_port, d(28) => 
                           from_mux_2_1_to_latch_high_28_port, d(27) => 
                           from_mux_2_1_to_latch_high_27_port, d(26) => 
                           from_mux_2_1_to_latch_high_26_port, d(25) => 
                           from_mux_2_1_to_latch_high_25_port, d(24) => 
                           from_mux_2_1_to_latch_high_24_port, d(23) => 
                           from_mux_2_1_to_latch_high_23_port, d(22) => 
                           from_mux_2_1_to_latch_high_22_port, d(21) => 
                           from_mux_2_1_to_latch_high_21_port, d(20) => 
                           from_mux_2_1_to_latch_high_20_port, d(19) => 
                           from_mux_2_1_to_latch_high_19_port, d(18) => 
                           from_mux_2_1_to_latch_high_18_port, d(17) => 
                           from_mux_2_1_to_latch_high_17_port, d(16) => 
                           from_mux_2_1_to_latch_high_16_port, d(15) => 
                           from_mux_2_1_to_latch_high_15_port, d(14) => 
                           from_mux_2_1_to_latch_high_14_port, d(13) => 
                           from_mux_2_1_to_latch_high_13_port, d(12) => 
                           from_mux_2_1_to_latch_high_12_port, d(11) => 
                           from_mux_2_1_to_latch_high_11_port, d(10) => 
                           from_mux_2_1_to_latch_high_10_port, d(9) => 
                           from_mux_2_1_to_latch_high_9_port, d(8) => 
                           from_mux_2_1_to_latch_high_8_port, d(7) => 
                           from_mux_2_1_to_latch_high_7_port, d(6) => 
                           from_mux_2_1_to_latch_high_6_port, d(5) => 
                           from_mux_2_1_to_latch_high_5_port, d(4) => 
                           from_mux_2_1_to_latch_high_4_port, d(3) => 
                           from_mux_2_1_to_latch_high_3_port, d(2) => 
                           from_mux_2_1_to_latch_high_2_port, d(1) => 
                           from_mux_2_1_to_latch_high_1_port, d(0) => 
                           from_mux_2_1_to_latch_high_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => net2756, q(30) => 
                           net2757, q(29) => net2758, q(28) => net2759, q(27) 
                           => net2760, q(26) => net2761, q(25) => net2762, 
                           q(24) => net2763, q(23) => net2764, q(22) => net2765
                           , q(21) => net2766, q(20) => net2767, q(19) => 
                           net2768, q(18) => net2769, q(17) => net2770, q(16) 
                           => net2771, q(15) => from_latch_to_mul_op1_15_port, 
                           q(14) => from_latch_to_mul_op1_14_port, q(13) => 
                           from_latch_to_mul_op1_13_port, q(12) => 
                           from_latch_to_mul_op1_12_port, q(11) => 
                           from_latch_to_mul_op1_11_port, q(10) => 
                           from_latch_to_mul_op1_10_port, q(9) => 
                           from_latch_to_mul_op1_9_port, q(8) => 
                           from_latch_to_mul_op1_8_port, q(7) => 
                           from_latch_to_mul_op1_7_port, q(6) => 
                           from_latch_to_mul_op1_6_port, q(5) => 
                           from_latch_to_mul_op1_5_port, q(4) => 
                           from_latch_to_mul_op1_4_port, q(3) => 
                           from_latch_to_mul_op1_3_port, q(2) => 
                           from_latch_to_mul_op1_2_port, q(1) => 
                           from_latch_to_mul_op1_1_port, q(0) => 
                           from_latch_to_mul_op1_0_port);
   PL5 : positive_latch_on_010_1 port map( d(31) => 
                           from_mux_2_1_to_latch_low_31_port, d(30) => 
                           from_mux_2_1_to_latch_low_30_port, d(29) => 
                           from_mux_2_1_to_latch_low_29_port, d(28) => 
                           from_mux_2_1_to_latch_low_28_port, d(27) => 
                           from_mux_2_1_to_latch_low_27_port, d(26) => 
                           from_mux_2_1_to_latch_low_26_port, d(25) => 
                           from_mux_2_1_to_latch_low_25_port, d(24) => 
                           from_mux_2_1_to_latch_low_24_port, d(23) => 
                           from_mux_2_1_to_latch_low_23_port, d(22) => 
                           from_mux_2_1_to_latch_low_22_port, d(21) => 
                           from_mux_2_1_to_latch_low_21_port, d(20) => 
                           from_mux_2_1_to_latch_low_20_port, d(19) => 
                           from_mux_2_1_to_latch_low_19_port, d(18) => 
                           from_mux_2_1_to_latch_low_18_port, d(17) => 
                           from_mux_2_1_to_latch_low_17_port, d(16) => 
                           from_mux_2_1_to_latch_low_16_port, d(15) => 
                           from_mux_2_1_to_latch_low_15_port, d(14) => 
                           from_mux_2_1_to_latch_low_14_port, d(13) => 
                           from_mux_2_1_to_latch_low_13_port, d(12) => 
                           from_mux_2_1_to_latch_low_12_port, d(11) => 
                           from_mux_2_1_to_latch_low_11_port, d(10) => 
                           from_mux_2_1_to_latch_low_10_port, d(9) => 
                           from_mux_2_1_to_latch_low_9_port, d(8) => 
                           from_mux_2_1_to_latch_low_8_port, d(7) => 
                           from_mux_2_1_to_latch_low_7_port, d(6) => 
                           from_mux_2_1_to_latch_low_6_port, d(5) => 
                           from_mux_2_1_to_latch_low_5_port, d(4) => 
                           from_mux_2_1_to_latch_low_4_port, d(3) => 
                           from_mux_2_1_to_latch_low_3_port, d(2) => 
                           from_mux_2_1_to_latch_low_2_port, d(1) => 
                           from_mux_2_1_to_latch_low_1_port, d(0) => 
                           from_mux_2_1_to_latch_low_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => net2740, q(30) => 
                           net2741, q(29) => net2742, q(28) => net2743, q(27) 
                           => net2744, q(26) => net2745, q(25) => net2746, 
                           q(24) => net2747, q(23) => net2748, q(22) => net2749
                           , q(21) => net2750, q(20) => net2751, q(19) => 
                           net2752, q(18) => net2753, q(17) => net2754, q(16) 
                           => net2755, q(15) => from_latch_to_mul_op2_15_port, 
                           q(14) => from_latch_to_mul_op2_14_port, q(13) => 
                           from_latch_to_mul_op2_13_port, q(12) => 
                           from_latch_to_mul_op2_12_port, q(11) => 
                           from_latch_to_mul_op2_11_port, q(10) => 
                           from_latch_to_mul_op2_10_port, q(9) => 
                           from_latch_to_mul_op2_9_port, q(8) => 
                           from_latch_to_mul_op2_8_port, q(7) => 
                           from_latch_to_mul_op2_7_port, q(6) => 
                           from_latch_to_mul_op2_6_port, q(5) => 
                           from_latch_to_mul_op2_5_port, q(4) => 
                           from_latch_to_mul_op2_4_port, q(3) => 
                           from_latch_to_mul_op2_3_port, q(2) => 
                           from_latch_to_mul_op2_2_port, q(1) => 
                           from_latch_to_mul_op2_1_port, q(0) => 
                           from_latch_to_mul_op2_0_port);
   PL6 : positive_latch_on_011_0 port map( d(31) => 
                           from_mux_2_1_to_latch_high_31_port, d(30) => 
                           from_mux_2_1_to_latch_high_30_port, d(29) => 
                           from_mux_2_1_to_latch_high_29_port, d(28) => 
                           from_mux_2_1_to_latch_high_28_port, d(27) => 
                           from_mux_2_1_to_latch_high_27_port, d(26) => 
                           from_mux_2_1_to_latch_high_26_port, d(25) => 
                           from_mux_2_1_to_latch_high_25_port, d(24) => 
                           from_mux_2_1_to_latch_high_24_port, d(23) => 
                           from_mux_2_1_to_latch_high_23_port, d(22) => 
                           from_mux_2_1_to_latch_high_22_port, d(21) => 
                           from_mux_2_1_to_latch_high_21_port, d(20) => 
                           from_mux_2_1_to_latch_high_20_port, d(19) => 
                           from_mux_2_1_to_latch_high_19_port, d(18) => 
                           from_mux_2_1_to_latch_high_18_port, d(17) => 
                           from_mux_2_1_to_latch_high_17_port, d(16) => 
                           from_mux_2_1_to_latch_high_16_port, d(15) => 
                           from_mux_2_1_to_latch_high_15_port, d(14) => 
                           from_mux_2_1_to_latch_high_14_port, d(13) => 
                           from_mux_2_1_to_latch_high_13_port, d(12) => 
                           from_mux_2_1_to_latch_high_12_port, d(11) => 
                           from_mux_2_1_to_latch_high_11_port, d(10) => 
                           from_mux_2_1_to_latch_high_10_port, d(9) => 
                           from_mux_2_1_to_latch_high_9_port, d(8) => 
                           from_mux_2_1_to_latch_high_8_port, d(7) => 
                           from_mux_2_1_to_latch_high_7_port, d(6) => 
                           from_mux_2_1_to_latch_high_6_port, d(5) => 
                           from_mux_2_1_to_latch_high_5_port, d(4) => 
                           from_mux_2_1_to_latch_high_4_port, d(3) => 
                           from_mux_2_1_to_latch_high_3_port, d(2) => 
                           from_mux_2_1_to_latch_high_2_port, d(1) => 
                           from_mux_2_1_to_latch_high_1_port, d(0) => 
                           from_mux_2_1_to_latch_high_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_shifter_op1_31_port, q(30) => 
                           from_latch_to_shifter_op1_30_port, q(29) => 
                           from_latch_to_shifter_op1_29_port, q(28) => 
                           from_latch_to_shifter_op1_28_port, q(27) => 
                           from_latch_to_shifter_op1_27_port, q(26) => 
                           from_latch_to_shifter_op1_26_port, q(25) => 
                           from_latch_to_shifter_op1_25_port, q(24) => 
                           from_latch_to_shifter_op1_24_port, q(23) => 
                           from_latch_to_shifter_op1_23_port, q(22) => 
                           from_latch_to_shifter_op1_22_port, q(21) => 
                           from_latch_to_shifter_op1_21_port, q(20) => 
                           from_latch_to_shifter_op1_20_port, q(19) => 
                           from_latch_to_shifter_op1_19_port, q(18) => 
                           from_latch_to_shifter_op1_18_port, q(17) => 
                           from_latch_to_shifter_op1_17_port, q(16) => 
                           from_latch_to_shifter_op1_16_port, q(15) => 
                           from_latch_to_shifter_op1_15_port, q(14) => 
                           from_latch_to_shifter_op1_14_port, q(13) => 
                           from_latch_to_shifter_op1_13_port, q(12) => 
                           from_latch_to_shifter_op1_12_port, q(11) => 
                           from_latch_to_shifter_op1_11_port, q(10) => 
                           from_latch_to_shifter_op1_10_port, q(9) => 
                           from_latch_to_shifter_op1_9_port, q(8) => 
                           from_latch_to_shifter_op1_8_port, q(7) => 
                           from_latch_to_shifter_op1_7_port, q(6) => 
                           from_latch_to_shifter_op1_6_port, q(5) => 
                           from_latch_to_shifter_op1_5_port, q(4) => 
                           from_latch_to_shifter_op1_4_port, q(3) => 
                           from_latch_to_shifter_op1_3_port, q(2) => 
                           from_latch_to_shifter_op1_2_port, q(1) => 
                           from_latch_to_shifter_op1_1_port, q(0) => 
                           from_latch_to_shifter_op1_0_port);
   PL7 : positive_latch_on_011_1 port map( d(31) => 
                           from_mux_2_1_to_latch_low_31_port, d(30) => 
                           from_mux_2_1_to_latch_low_30_port, d(29) => 
                           from_mux_2_1_to_latch_low_29_port, d(28) => 
                           from_mux_2_1_to_latch_low_28_port, d(27) => 
                           from_mux_2_1_to_latch_low_27_port, d(26) => 
                           from_mux_2_1_to_latch_low_26_port, d(25) => 
                           from_mux_2_1_to_latch_low_25_port, d(24) => 
                           from_mux_2_1_to_latch_low_24_port, d(23) => 
                           from_mux_2_1_to_latch_low_23_port, d(22) => 
                           from_mux_2_1_to_latch_low_22_port, d(21) => 
                           from_mux_2_1_to_latch_low_21_port, d(20) => 
                           from_mux_2_1_to_latch_low_20_port, d(19) => 
                           from_mux_2_1_to_latch_low_19_port, d(18) => 
                           from_mux_2_1_to_latch_low_18_port, d(17) => 
                           from_mux_2_1_to_latch_low_17_port, d(16) => 
                           from_mux_2_1_to_latch_low_16_port, d(15) => 
                           from_mux_2_1_to_latch_low_15_port, d(14) => 
                           from_mux_2_1_to_latch_low_14_port, d(13) => 
                           from_mux_2_1_to_latch_low_13_port, d(12) => 
                           from_mux_2_1_to_latch_low_12_port, d(11) => 
                           from_mux_2_1_to_latch_low_11_port, d(10) => 
                           from_mux_2_1_to_latch_low_10_port, d(9) => 
                           from_mux_2_1_to_latch_low_9_port, d(8) => 
                           from_mux_2_1_to_latch_low_8_port, d(7) => 
                           from_mux_2_1_to_latch_low_7_port, d(6) => 
                           from_mux_2_1_to_latch_low_6_port, d(5) => 
                           from_mux_2_1_to_latch_low_5_port, d(4) => 
                           from_mux_2_1_to_latch_low_4_port, d(3) => 
                           from_mux_2_1_to_latch_low_3_port, d(2) => 
                           from_mux_2_1_to_latch_low_2_port, d(1) => 
                           from_mux_2_1_to_latch_low_1_port, d(0) => 
                           from_mux_2_1_to_latch_low_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_shifter_op2_31_port, q(30) => 
                           from_latch_to_shifter_op2_30_port, q(29) => 
                           from_latch_to_shifter_op2_29_port, q(28) => 
                           from_latch_to_shifter_op2_28_port, q(27) => 
                           from_latch_to_shifter_op2_27_port, q(26) => 
                           from_latch_to_shifter_op2_26_port, q(25) => 
                           from_latch_to_shifter_op2_25_port, q(24) => 
                           from_latch_to_shifter_op2_24_port, q(23) => 
                           from_latch_to_shifter_op2_23_port, q(22) => 
                           from_latch_to_shifter_op2_22_port, q(21) => 
                           from_latch_to_shifter_op2_21_port, q(20) => 
                           from_latch_to_shifter_op2_20_port, q(19) => 
                           from_latch_to_shifter_op2_19_port, q(18) => 
                           from_latch_to_shifter_op2_18_port, q(17) => 
                           from_latch_to_shifter_op2_17_port, q(16) => 
                           from_latch_to_shifter_op2_16_port, q(15) => 
                           from_latch_to_shifter_op2_15_port, q(14) => 
                           from_latch_to_shifter_op2_14_port, q(13) => 
                           from_latch_to_shifter_op2_13_port, q(12) => 
                           from_latch_to_shifter_op2_12_port, q(11) => 
                           from_latch_to_shifter_op2_11_port, q(10) => 
                           from_latch_to_shifter_op2_10_port, q(9) => 
                           from_latch_to_shifter_op2_9_port, q(8) => 
                           from_latch_to_shifter_op2_8_port, q(7) => 
                           from_latch_to_shifter_op2_7_port, q(6) => 
                           from_latch_to_shifter_op2_6_port, q(5) => 
                           from_latch_to_shifter_op2_5_port, q(4) => 
                           from_latch_to_shifter_op2_4_port, q(3) => 
                           from_latch_to_shifter_op2_3_port, q(2) => 
                           from_latch_to_shifter_op2_2_port, q(1) => 
                           from_latch_to_shifter_op2_1_port, q(0) => 
                           from_latch_to_shifter_op2_0_port);
   PL8 : positive_latch_on_100_0 port map( d(31) => 
                           from_mux_2_1_to_latch_high_31_port, d(30) => 
                           from_mux_2_1_to_latch_high_30_port, d(29) => 
                           from_mux_2_1_to_latch_high_29_port, d(28) => 
                           from_mux_2_1_to_latch_high_28_port, d(27) => 
                           from_mux_2_1_to_latch_high_27_port, d(26) => 
                           from_mux_2_1_to_latch_high_26_port, d(25) => 
                           from_mux_2_1_to_latch_high_25_port, d(24) => 
                           from_mux_2_1_to_latch_high_24_port, d(23) => 
                           from_mux_2_1_to_latch_high_23_port, d(22) => 
                           from_mux_2_1_to_latch_high_22_port, d(21) => 
                           from_mux_2_1_to_latch_high_21_port, d(20) => 
                           from_mux_2_1_to_latch_high_20_port, d(19) => 
                           from_mux_2_1_to_latch_high_19_port, d(18) => 
                           from_mux_2_1_to_latch_high_18_port, d(17) => 
                           from_mux_2_1_to_latch_high_17_port, d(16) => 
                           from_mux_2_1_to_latch_high_16_port, d(15) => 
                           from_mux_2_1_to_latch_high_15_port, d(14) => 
                           from_mux_2_1_to_latch_high_14_port, d(13) => 
                           from_mux_2_1_to_latch_high_13_port, d(12) => 
                           from_mux_2_1_to_latch_high_12_port, d(11) => 
                           from_mux_2_1_to_latch_high_11_port, d(10) => 
                           from_mux_2_1_to_latch_high_10_port, d(9) => 
                           from_mux_2_1_to_latch_high_9_port, d(8) => 
                           from_mux_2_1_to_latch_high_8_port, d(7) => 
                           from_mux_2_1_to_latch_high_7_port, d(6) => 
                           from_mux_2_1_to_latch_high_6_port, d(5) => 
                           from_mux_2_1_to_latch_high_5_port, d(4) => 
                           from_mux_2_1_to_latch_high_4_port, d(3) => 
                           from_mux_2_1_to_latch_high_3_port, d(2) => 
                           from_mux_2_1_to_latch_high_2_port, d(1) => 
                           from_mux_2_1_to_latch_high_1_port, d(0) => 
                           from_mux_2_1_to_latch_high_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_comparator_op1_31_port, q(30) => 
                           from_latch_to_comparator_op1_30_port, q(29) => 
                           from_latch_to_comparator_op1_29_port, q(28) => 
                           from_latch_to_comparator_op1_28_port, q(27) => 
                           from_latch_to_comparator_op1_27_port, q(26) => 
                           from_latch_to_comparator_op1_26_port, q(25) => 
                           from_latch_to_comparator_op1_25_port, q(24) => 
                           from_latch_to_comparator_op1_24_port, q(23) => 
                           from_latch_to_comparator_op1_23_port, q(22) => 
                           from_latch_to_comparator_op1_22_port, q(21) => 
                           from_latch_to_comparator_op1_21_port, q(20) => 
                           from_latch_to_comparator_op1_20_port, q(19) => 
                           from_latch_to_comparator_op1_19_port, q(18) => 
                           from_latch_to_comparator_op1_18_port, q(17) => 
                           from_latch_to_comparator_op1_17_port, q(16) => 
                           from_latch_to_comparator_op1_16_port, q(15) => 
                           from_latch_to_comparator_op1_15_port, q(14) => 
                           from_latch_to_comparator_op1_14_port, q(13) => 
                           from_latch_to_comparator_op1_13_port, q(12) => 
                           from_latch_to_comparator_op1_12_port, q(11) => 
                           from_latch_to_comparator_op1_11_port, q(10) => 
                           from_latch_to_comparator_op1_10_port, q(9) => 
                           from_latch_to_comparator_op1_9_port, q(8) => 
                           from_latch_to_comparator_op1_8_port, q(7) => 
                           from_latch_to_comparator_op1_7_port, q(6) => 
                           from_latch_to_comparator_op1_6_port, q(5) => 
                           from_latch_to_comparator_op1_5_port, q(4) => 
                           from_latch_to_comparator_op1_4_port, q(3) => 
                           from_latch_to_comparator_op1_3_port, q(2) => 
                           from_latch_to_comparator_op1_2_port, q(1) => 
                           from_latch_to_comparator_op1_1_port, q(0) => 
                           from_latch_to_comparator_op1_0_port);
   PL9 : positive_latch_on_100_1 port map( d(31) => 
                           from_mux_2_1_to_latch_low_31_port, d(30) => 
                           from_mux_2_1_to_latch_low_30_port, d(29) => 
                           from_mux_2_1_to_latch_low_29_port, d(28) => 
                           from_mux_2_1_to_latch_low_28_port, d(27) => 
                           from_mux_2_1_to_latch_low_27_port, d(26) => 
                           from_mux_2_1_to_latch_low_26_port, d(25) => 
                           from_mux_2_1_to_latch_low_25_port, d(24) => 
                           from_mux_2_1_to_latch_low_24_port, d(23) => 
                           from_mux_2_1_to_latch_low_23_port, d(22) => 
                           from_mux_2_1_to_latch_low_22_port, d(21) => 
                           from_mux_2_1_to_latch_low_21_port, d(20) => 
                           from_mux_2_1_to_latch_low_20_port, d(19) => 
                           from_mux_2_1_to_latch_low_19_port, d(18) => 
                           from_mux_2_1_to_latch_low_18_port, d(17) => 
                           from_mux_2_1_to_latch_low_17_port, d(16) => 
                           from_mux_2_1_to_latch_low_16_port, d(15) => 
                           from_mux_2_1_to_latch_low_15_port, d(14) => 
                           from_mux_2_1_to_latch_low_14_port, d(13) => 
                           from_mux_2_1_to_latch_low_13_port, d(12) => 
                           from_mux_2_1_to_latch_low_12_port, d(11) => 
                           from_mux_2_1_to_latch_low_11_port, d(10) => 
                           from_mux_2_1_to_latch_low_10_port, d(9) => 
                           from_mux_2_1_to_latch_low_9_port, d(8) => 
                           from_mux_2_1_to_latch_low_8_port, d(7) => 
                           from_mux_2_1_to_latch_low_7_port, d(6) => 
                           from_mux_2_1_to_latch_low_6_port, d(5) => 
                           from_mux_2_1_to_latch_low_5_port, d(4) => 
                           from_mux_2_1_to_latch_low_4_port, d(3) => 
                           from_mux_2_1_to_latch_low_3_port, d(2) => 
                           from_mux_2_1_to_latch_low_2_port, d(1) => 
                           from_mux_2_1_to_latch_low_1_port, d(0) => 
                           from_mux_2_1_to_latch_low_0_port, enable(2) => 
                           sel_signal_5_1_2_port, enable(1) => 
                           sel_signal_5_1_1_port, enable(0) => 
                           sel_signal_5_1_0_port, q(31) => 
                           from_latch_to_comparator_op2_31_port, q(30) => 
                           from_latch_to_comparator_op2_30_port, q(29) => 
                           from_latch_to_comparator_op2_29_port, q(28) => 
                           from_latch_to_comparator_op2_28_port, q(27) => 
                           from_latch_to_comparator_op2_27_port, q(26) => 
                           from_latch_to_comparator_op2_26_port, q(25) => 
                           from_latch_to_comparator_op2_25_port, q(24) => 
                           from_latch_to_comparator_op2_24_port, q(23) => 
                           from_latch_to_comparator_op2_23_port, q(22) => 
                           from_latch_to_comparator_op2_22_port, q(21) => 
                           from_latch_to_comparator_op2_21_port, q(20) => 
                           from_latch_to_comparator_op2_20_port, q(19) => 
                           from_latch_to_comparator_op2_19_port, q(18) => 
                           from_latch_to_comparator_op2_18_port, q(17) => 
                           from_latch_to_comparator_op2_17_port, q(16) => 
                           from_latch_to_comparator_op2_16_port, q(15) => 
                           from_latch_to_comparator_op2_15_port, q(14) => 
                           from_latch_to_comparator_op2_14_port, q(13) => 
                           from_latch_to_comparator_op2_13_port, q(12) => 
                           from_latch_to_comparator_op2_12_port, q(11) => 
                           from_latch_to_comparator_op2_11_port, q(10) => 
                           from_latch_to_comparator_op2_10_port, q(9) => 
                           from_latch_to_comparator_op2_9_port, q(8) => 
                           from_latch_to_comparator_op2_8_port, q(7) => 
                           from_latch_to_comparator_op2_7_port, q(6) => 
                           from_latch_to_comparator_op2_6_port, q(5) => 
                           from_latch_to_comparator_op2_5_port, q(4) => 
                           from_latch_to_comparator_op2_4_port, q(3) => 
                           from_latch_to_comparator_op2_3_port, q(2) => 
                           from_latch_to_comparator_op2_2_port, q(1) => 
                           from_latch_to_comparator_op2_1_port, q(0) => 
                           from_latch_to_comparator_op2_0_port);
   COMP : comparator port map( A(31) => from_latch_to_comparator_op1_31_port, 
                           A(30) => from_latch_to_comparator_op1_30_port, A(29)
                           => from_latch_to_comparator_op1_29_port, A(28) => 
                           from_latch_to_comparator_op1_28_port, A(27) => 
                           from_latch_to_comparator_op1_27_port, A(26) => 
                           from_latch_to_comparator_op1_26_port, A(25) => 
                           from_latch_to_comparator_op1_25_port, A(24) => 
                           from_latch_to_comparator_op1_24_port, A(23) => 
                           from_latch_to_comparator_op1_23_port, A(22) => 
                           from_latch_to_comparator_op1_22_port, A(21) => 
                           from_latch_to_comparator_op1_21_port, A(20) => 
                           from_latch_to_comparator_op1_20_port, A(19) => 
                           from_latch_to_comparator_op1_19_port, A(18) => 
                           from_latch_to_comparator_op1_18_port, A(17) => 
                           from_latch_to_comparator_op1_17_port, A(16) => 
                           from_latch_to_comparator_op1_16_port, A(15) => 
                           from_latch_to_comparator_op1_15_port, A(14) => 
                           from_latch_to_comparator_op1_14_port, A(13) => 
                           from_latch_to_comparator_op1_13_port, A(12) => 
                           from_latch_to_comparator_op1_12_port, A(11) => 
                           from_latch_to_comparator_op1_11_port, A(10) => 
                           from_latch_to_comparator_op1_10_port, A(9) => 
                           from_latch_to_comparator_op1_9_port, A(8) => 
                           from_latch_to_comparator_op1_8_port, A(7) => 
                           from_latch_to_comparator_op1_7_port, A(6) => 
                           from_latch_to_comparator_op1_6_port, A(5) => 
                           from_latch_to_comparator_op1_5_port, A(4) => 
                           from_latch_to_comparator_op1_4_port, A(3) => 
                           from_latch_to_comparator_op1_3_port, A(2) => 
                           from_latch_to_comparator_op1_2_port, A(1) => 
                           from_latch_to_comparator_op1_1_port, A(0) => 
                           from_latch_to_comparator_op1_0_port, B(31) => 
                           from_latch_to_comparator_op2_31_port, B(30) => 
                           from_latch_to_comparator_op2_30_port, B(29) => 
                           from_latch_to_comparator_op2_29_port, B(28) => 
                           from_latch_to_comparator_op2_28_port, B(27) => 
                           from_latch_to_comparator_op2_27_port, B(26) => 
                           from_latch_to_comparator_op2_26_port, B(25) => 
                           from_latch_to_comparator_op2_25_port, B(24) => 
                           from_latch_to_comparator_op2_24_port, B(23) => 
                           from_latch_to_comparator_op2_23_port, B(22) => 
                           from_latch_to_comparator_op2_22_port, B(21) => 
                           from_latch_to_comparator_op2_21_port, B(20) => 
                           from_latch_to_comparator_op2_20_port, B(19) => 
                           from_latch_to_comparator_op2_19_port, B(18) => 
                           from_latch_to_comparator_op2_18_port, B(17) => 
                           from_latch_to_comparator_op2_17_port, B(16) => 
                           from_latch_to_comparator_op2_16_port, B(15) => 
                           from_latch_to_comparator_op2_15_port, B(14) => 
                           from_latch_to_comparator_op2_14_port, B(13) => 
                           from_latch_to_comparator_op2_13_port, B(12) => 
                           from_latch_to_comparator_op2_12_port, B(11) => 
                           from_latch_to_comparator_op2_11_port, B(10) => 
                           from_latch_to_comparator_op2_10_port, B(9) => 
                           from_latch_to_comparator_op2_9_port, B(8) => 
                           from_latch_to_comparator_op2_8_port, B(7) => 
                           from_latch_to_comparator_op2_7_port, B(6) => 
                           from_latch_to_comparator_op2_6_port, B(5) => 
                           from_latch_to_comparator_op2_5_port, B(4) => 
                           from_latch_to_comparator_op2_4_port, B(3) => 
                           from_latch_to_comparator_op2_3_port, B(2) => 
                           from_latch_to_comparator_op2_2_port, B(1) => 
                           from_latch_to_comparator_op2_1_port, B(0) => 
                           from_latch_to_comparator_op2_0_port, Sel(2) => 
                           sel_comparator_2_port, Sel(1) => 
                           sel_comparator_1_port, Sel(0) => 
                           sel_comparator_0_port, O(31) => n_1056, O(30) => 
                           n_1057, O(29) => n_1058, O(28) => n_1059, O(27) => 
                           n_1060, O(26) => n_1061, O(25) => n_1062, O(24) => 
                           n_1063, O(23) => n_1064, O(22) => n_1065, O(21) => 
                           n_1066, O(20) => n_1067, O(19) => n_1068, O(18) => 
                           n_1069, O(17) => n_1070, O(16) => n_1071, O(15) => 
                           n_1072, O(14) => n_1073, O(13) => n_1074, O(12) => 
                           n_1075, O(11) => n_1076, O(10) => n_1077, O(9) => 
                           n_1078, O(8) => n_1079, O(7) => n_1080, O(6) => 
                           n_1081, O(5) => n_1082, O(4) => n_1083, O(3) => 
                           n_1084, O(2) => n_1085, O(1) => n_1086, O(0) => 
                           jump_port);
   P4 : pentium4_adder_XBIT32_NBIT4_0 port map( A(31) => 
                           from_latch_to_adder_op1_31_port, A(30) => 
                           from_latch_to_adder_op1_30_port, A(29) => 
                           from_latch_to_adder_op1_29_port, A(28) => 
                           from_latch_to_adder_op1_28_port, A(27) => 
                           from_latch_to_adder_op1_27_port, A(26) => 
                           from_latch_to_adder_op1_26_port, A(25) => 
                           from_latch_to_adder_op1_25_port, A(24) => 
                           from_latch_to_adder_op1_24_port, A(23) => 
                           from_latch_to_adder_op1_23_port, A(22) => 
                           from_latch_to_adder_op1_22_port, A(21) => 
                           from_latch_to_adder_op1_21_port, A(20) => 
                           from_latch_to_adder_op1_20_port, A(19) => 
                           from_latch_to_adder_op1_19_port, A(18) => 
                           from_latch_to_adder_op1_18_port, A(17) => 
                           from_latch_to_adder_op1_17_port, A(16) => 
                           from_latch_to_adder_op1_16_port, A(15) => 
                           from_latch_to_adder_op1_15_port, A(14) => 
                           from_latch_to_adder_op1_14_port, A(13) => 
                           from_latch_to_adder_op1_13_port, A(12) => 
                           from_latch_to_adder_op1_12_port, A(11) => 
                           from_latch_to_adder_op1_11_port, A(10) => 
                           from_latch_to_adder_op1_10_port, A(9) => 
                           from_latch_to_adder_op1_9_port, A(8) => 
                           from_latch_to_adder_op1_8_port, A(7) => 
                           from_latch_to_adder_op1_7_port, A(6) => 
                           from_latch_to_adder_op1_6_port, A(5) => 
                           from_latch_to_adder_op1_5_port, A(4) => 
                           from_latch_to_adder_op1_4_port, A(3) => 
                           from_latch_to_adder_op1_3_port, A(2) => 
                           from_latch_to_adder_op1_2_port, A(1) => 
                           from_latch_to_adder_op1_1_port, A(0) => 
                           from_latch_to_adder_op1_0_port, B(31) => 
                           from_latch_to_mux_sub_or_add_31_port, B(30) => 
                           from_latch_to_mux_sub_or_add_30_port, B(29) => 
                           from_latch_to_mux_sub_or_add_29_port, B(28) => 
                           from_latch_to_mux_sub_or_add_28_port, B(27) => 
                           from_latch_to_mux_sub_or_add_27_port, B(26) => 
                           from_latch_to_mux_sub_or_add_26_port, B(25) => 
                           from_latch_to_mux_sub_or_add_25_port, B(24) => 
                           from_latch_to_mux_sub_or_add_24_port, B(23) => 
                           from_latch_to_mux_sub_or_add_23_port, B(22) => 
                           from_latch_to_mux_sub_or_add_22_port, B(21) => 
                           from_latch_to_mux_sub_or_add_21_port, B(20) => 
                           from_latch_to_mux_sub_or_add_20_port, B(19) => 
                           from_latch_to_mux_sub_or_add_19_port, B(18) => 
                           from_latch_to_mux_sub_or_add_18_port, B(17) => 
                           from_latch_to_mux_sub_or_add_17_port, B(16) => 
                           from_latch_to_mux_sub_or_add_16_port, B(15) => 
                           from_latch_to_mux_sub_or_add_15_port, B(14) => 
                           from_latch_to_mux_sub_or_add_14_port, B(13) => 
                           from_latch_to_mux_sub_or_add_13_port, B(12) => 
                           from_latch_to_mux_sub_or_add_12_port, B(11) => 
                           from_latch_to_mux_sub_or_add_11_port, B(10) => 
                           from_latch_to_mux_sub_or_add_10_port, B(9) => 
                           from_latch_to_mux_sub_or_add_9_port, B(8) => 
                           from_latch_to_mux_sub_or_add_8_port, B(7) => 
                           from_latch_to_mux_sub_or_add_7_port, B(6) => 
                           from_latch_to_mux_sub_or_add_6_port, B(5) => 
                           from_latch_to_mux_sub_or_add_5_port, B(4) => 
                           from_latch_to_mux_sub_or_add_4_port, B(3) => 
                           from_latch_to_mux_sub_or_add_3_port, B(2) => 
                           from_latch_to_mux_sub_or_add_2_port, B(1) => 
                           from_latch_to_mux_sub_or_add_1_port, B(0) => 
                           from_latch_to_mux_sub_or_add_0_port, C_0 => carry_in
                           , S(31) => from_adder_to_mux_31_port, S(30) => 
                           from_adder_to_mux_30_port, S(29) => 
                           from_adder_to_mux_29_port, S(28) => 
                           from_adder_to_mux_28_port, S(27) => 
                           from_adder_to_mux_27_port, S(26) => 
                           from_adder_to_mux_26_port, S(25) => 
                           from_adder_to_mux_25_port, S(24) => 
                           from_adder_to_mux_24_port, S(23) => 
                           from_adder_to_mux_23_port, S(22) => 
                           from_adder_to_mux_22_port, S(21) => 
                           from_adder_to_mux_21_port, S(20) => 
                           from_adder_to_mux_20_port, S(19) => 
                           from_adder_to_mux_19_port, S(18) => 
                           from_adder_to_mux_18_port, S(17) => 
                           from_adder_to_mux_17_port, S(16) => 
                           from_adder_to_mux_16_port, S(15) => 
                           from_adder_to_mux_15_port, S(14) => 
                           from_adder_to_mux_14_port, S(13) => 
                           from_adder_to_mux_13_port, S(12) => 
                           from_adder_to_mux_12_port, S(11) => 
                           from_adder_to_mux_11_port, S(10) => 
                           from_adder_to_mux_10_port, S(9) => 
                           from_adder_to_mux_9_port, S(8) => 
                           from_adder_to_mux_8_port, S(7) => 
                           from_adder_to_mux_7_port, S(6) => 
                           from_adder_to_mux_6_port, S(5) => 
                           from_adder_to_mux_5_port, S(4) => 
                           from_adder_to_mux_4_port, S(3) => 
                           from_adder_to_mux_3_port, S(2) => 
                           from_adder_to_mux_2_port, S(1) => 
                           from_adder_to_mux_1_port, S(0) => 
                           from_adder_to_mux_0_port, Cout => net2739);
   BRANCH_ADDER : pentium4_adder_XBIT32_NBIT4_8 port map( A(31) => 
                           operand_pc(31), A(30) => operand_pc(30), A(29) => 
                           operand_pc(29), A(28) => operand_pc(28), A(27) => 
                           operand_pc(27), A(26) => operand_pc(26), A(25) => 
                           operand_pc(25), A(24) => operand_pc(24), A(23) => 
                           operand_pc(23), A(22) => operand_pc(22), A(21) => 
                           operand_pc(21), A(20) => operand_pc(20), A(19) => 
                           operand_pc(19), A(18) => operand_pc(18), A(17) => 
                           operand_pc(17), A(16) => operand_pc(16), A(15) => 
                           operand_pc(15), A(14) => operand_pc(14), A(13) => 
                           operand_pc(13), A(12) => operand_pc(12), A(11) => 
                           operand_pc(11), A(10) => operand_pc(10), A(9) => 
                           operand_pc(9), A(8) => operand_pc(8), A(7) => 
                           operand_pc(7), A(6) => operand_pc(6), A(5) => 
                           operand_pc(5), A(4) => operand_pc(4), A(3) => 
                           operand_pc(3), A(2) => operand_pc(2), A(1) => 
                           operand_pc(1), A(0) => operand_pc(0), B(31) => 
                           operand_imm(31), B(30) => operand_imm(31), B(29) => 
                           operand_imm(31), B(28) => operand_imm(30), B(27) => 
                           operand_imm(29), B(26) => operand_imm(28), B(25) => 
                           operand_imm(27), B(24) => operand_imm(26), B(23) => 
                           operand_imm(25), B(22) => operand_imm(24), B(21) => 
                           operand_imm(23), B(20) => operand_imm(22), B(19) => 
                           operand_imm(21), B(18) => operand_imm(20), B(17) => 
                           operand_imm(19), B(16) => operand_imm(18), B(15) => 
                           operand_imm(17), B(14) => operand_imm(16), B(13) => 
                           operand_imm(15), B(12) => operand_imm(14), B(11) => 
                           operand_imm(13), B(10) => operand_imm(12), B(9) => 
                           operand_imm(11), B(8) => operand_imm(10), B(7) => 
                           operand_imm(9), B(6) => operand_imm(8), B(5) => 
                           operand_imm(7), B(4) => operand_imm(6), B(3) => 
                           operand_imm(5), B(2) => operand_imm(4), B(1) => 
                           operand_imm(3), B(0) => operand_imm(2), C_0 => n4, 
                           S(31) => next_pc(31), S(30) => next_pc(30), S(29) =>
                           next_pc(29), S(28) => next_pc(28), S(27) => 
                           next_pc(27), S(26) => next_pc(26), S(25) => 
                           next_pc(25), S(24) => next_pc(24), S(23) => 
                           next_pc(23), S(22) => next_pc(22), S(21) => 
                           next_pc(21), S(20) => next_pc(20), S(19) => 
                           next_pc(19), S(18) => next_pc(18), S(17) => 
                           next_pc(17), S(16) => next_pc(16), S(15) => 
                           next_pc(15), S(14) => next_pc(14), S(13) => 
                           next_pc(13), S(12) => next_pc(12), S(11) => 
                           next_pc(11), S(10) => next_pc(10), S(9) => 
                           next_pc(9), S(8) => next_pc(8), S(7) => next_pc(7), 
                           S(6) => next_pc(6), S(5) => next_pc(5), S(4) => 
                           next_pc(4), S(3) => next_pc(3), S(2) => next_pc(2), 
                           S(1) => next_pc(1), S(0) => next_pc(0), Cout => 
                           net2738);
   M2 : Mux2X1_4 port map( a(31) => mux_to_mux_high_31_port, a(30) => 
                           mux_to_mux_high_30_port, a(29) => 
                           mux_to_mux_high_29_port, a(28) => 
                           mux_to_mux_high_28_port, a(27) => 
                           mux_to_mux_high_27_port, a(26) => 
                           mux_to_mux_high_26_port, a(25) => 
                           mux_to_mux_high_25_port, a(24) => 
                           mux_to_mux_high_24_port, a(23) => 
                           mux_to_mux_high_23_port, a(22) => 
                           mux_to_mux_high_22_port, a(21) => 
                           mux_to_mux_high_21_port, a(20) => 
                           mux_to_mux_high_20_port, a(19) => 
                           mux_to_mux_high_19_port, a(18) => 
                           mux_to_mux_high_18_port, a(17) => 
                           mux_to_mux_high_17_port, a(16) => 
                           mux_to_mux_high_16_port, a(15) => 
                           mux_to_mux_high_15_port, a(14) => 
                           mux_to_mux_high_14_port, a(13) => 
                           mux_to_mux_high_13_port, a(12) => 
                           mux_to_mux_high_12_port, a(11) => 
                           mux_to_mux_high_11_port, a(10) => 
                           mux_to_mux_high_10_port, a(9) => 
                           mux_to_mux_high_9_port, a(8) => 
                           mux_to_mux_high_8_port, a(7) => 
                           mux_to_mux_high_7_port, a(6) => 
                           mux_to_mux_high_6_port, a(5) => 
                           mux_to_mux_high_5_port, a(4) => 
                           mux_to_mux_high_4_port, a(3) => 
                           mux_to_mux_high_3_port, a(2) => 
                           mux_to_mux_high_2_port, a(1) => 
                           mux_to_mux_high_1_port, a(0) => 
                           mux_to_mux_high_0_port, b(31) => operand_pc(31), 
                           b(30) => operand_pc(30), b(29) => operand_pc(29), 
                           b(28) => operand_pc(28), b(27) => operand_pc(27), 
                           b(26) => operand_pc(26), b(25) => operand_pc(25), 
                           b(24) => operand_pc(24), b(23) => operand_pc(23), 
                           b(22) => operand_pc(22), b(21) => operand_pc(21), 
                           b(20) => operand_pc(20), b(19) => operand_pc(19), 
                           b(18) => operand_pc(18), b(17) => operand_pc(17), 
                           b(16) => operand_pc(16), b(15) => operand_pc(15), 
                           b(14) => operand_pc(14), b(13) => operand_pc(13), 
                           b(12) => operand_pc(12), b(11) => operand_pc(11), 
                           b(10) => operand_pc(10), b(9) => operand_pc(9), b(8)
                           => operand_pc(8), b(7) => operand_pc(7), b(6) => 
                           operand_pc(6), b(5) => operand_pc(5), b(4) => 
                           operand_pc(4), b(3) => operand_pc(3), b(2) => 
                           operand_pc(2), b(1) => operand_pc(1), b(0) => 
                           operand_pc(0), sel => sel_1, o(31) => 
                           from_mux_2_1_to_latch_high_31_port, o(30) => 
                           from_mux_2_1_to_latch_high_30_port, o(29) => 
                           from_mux_2_1_to_latch_high_29_port, o(28) => 
                           from_mux_2_1_to_latch_high_28_port, o(27) => 
                           from_mux_2_1_to_latch_high_27_port, o(26) => 
                           from_mux_2_1_to_latch_high_26_port, o(25) => 
                           from_mux_2_1_to_latch_high_25_port, o(24) => 
                           from_mux_2_1_to_latch_high_24_port, o(23) => 
                           from_mux_2_1_to_latch_high_23_port, o(22) => 
                           from_mux_2_1_to_latch_high_22_port, o(21) => 
                           from_mux_2_1_to_latch_high_21_port, o(20) => 
                           from_mux_2_1_to_latch_high_20_port, o(19) => 
                           from_mux_2_1_to_latch_high_19_port, o(18) => 
                           from_mux_2_1_to_latch_high_18_port, o(17) => 
                           from_mux_2_1_to_latch_high_17_port, o(16) => 
                           from_mux_2_1_to_latch_high_16_port, o(15) => 
                           from_mux_2_1_to_latch_high_15_port, o(14) => 
                           from_mux_2_1_to_latch_high_14_port, o(13) => 
                           from_mux_2_1_to_latch_high_13_port, o(12) => 
                           from_mux_2_1_to_latch_high_12_port, o(11) => 
                           from_mux_2_1_to_latch_high_11_port, o(10) => 
                           from_mux_2_1_to_latch_high_10_port, o(9) => 
                           from_mux_2_1_to_latch_high_9_port, o(8) => 
                           from_mux_2_1_to_latch_high_8_port, o(7) => 
                           from_mux_2_1_to_latch_high_7_port, o(6) => 
                           from_mux_2_1_to_latch_high_6_port, o(5) => 
                           from_mux_2_1_to_latch_high_5_port, o(4) => 
                           from_mux_2_1_to_latch_high_4_port, o(3) => 
                           from_mux_2_1_to_latch_high_3_port, o(2) => 
                           from_mux_2_1_to_latch_high_2_port, o(1) => 
                           from_mux_2_1_to_latch_high_1_port, o(0) => 
                           from_mux_2_1_to_latch_high_0_port);
   M3 : Mux2X1_3 port map( a(31) => mux_to_mux_low_31_port, a(30) => 
                           mux_to_mux_low_30_port, a(29) => 
                           mux_to_mux_low_29_port, a(28) => 
                           mux_to_mux_low_28_port, a(27) => 
                           mux_to_mux_low_27_port, a(26) => 
                           mux_to_mux_low_26_port, a(25) => 
                           mux_to_mux_low_25_port, a(24) => 
                           mux_to_mux_low_24_port, a(23) => 
                           mux_to_mux_low_23_port, a(22) => 
                           mux_to_mux_low_22_port, a(21) => 
                           mux_to_mux_low_21_port, a(20) => 
                           mux_to_mux_low_20_port, a(19) => 
                           mux_to_mux_low_19_port, a(18) => 
                           mux_to_mux_low_18_port, a(17) => 
                           mux_to_mux_low_17_port, a(16) => 
                           mux_to_mux_low_16_port, a(15) => 
                           mux_to_mux_low_15_port, a(14) => 
                           mux_to_mux_low_14_port, a(13) => 
                           mux_to_mux_low_13_port, a(12) => 
                           mux_to_mux_low_12_port, a(11) => 
                           mux_to_mux_low_11_port, a(10) => 
                           mux_to_mux_low_10_port, a(9) => 
                           mux_to_mux_low_9_port, a(8) => mux_to_mux_low_8_port
                           , a(7) => mux_to_mux_low_7_port, a(6) => 
                           mux_to_mux_low_6_port, a(5) => mux_to_mux_low_5_port
                           , a(4) => mux_to_mux_low_4_port, a(3) => 
                           mux_to_mux_low_3_port, a(2) => mux_to_mux_low_2_port
                           , a(1) => mux_to_mux_low_1_port, a(0) => 
                           mux_to_mux_low_0_port, b(31) => operand_imm(31), 
                           b(30) => operand_imm(30), b(29) => operand_imm(29), 
                           b(28) => operand_imm(28), b(27) => operand_imm(27), 
                           b(26) => operand_imm(26), b(25) => operand_imm(25), 
                           b(24) => operand_imm(24), b(23) => operand_imm(23), 
                           b(22) => operand_imm(22), b(21) => operand_imm(21), 
                           b(20) => operand_imm(20), b(19) => operand_imm(19), 
                           b(18) => operand_imm(18), b(17) => operand_imm(17), 
                           b(16) => operand_imm(16), b(15) => operand_imm(15), 
                           b(14) => operand_imm(14), b(13) => operand_imm(13), 
                           b(12) => operand_imm(12), b(11) => operand_imm(11), 
                           b(10) => operand_imm(10), b(9) => operand_imm(9), 
                           b(8) => operand_imm(8), b(7) => operand_imm(7), b(6)
                           => operand_imm(6), b(5) => operand_imm(5), b(4) => 
                           operand_imm(4), b(3) => operand_imm(3), b(2) => 
                           operand_imm(2), b(1) => operand_imm(1), b(0) => 
                           operand_imm(0), sel => sel_2, o(31) => 
                           from_mux_2_1_to_latch_low_31_port, o(30) => 
                           from_mux_2_1_to_latch_low_30_port, o(29) => 
                           from_mux_2_1_to_latch_low_29_port, o(28) => 
                           from_mux_2_1_to_latch_low_28_port, o(27) => 
                           from_mux_2_1_to_latch_low_27_port, o(26) => 
                           from_mux_2_1_to_latch_low_26_port, o(25) => 
                           from_mux_2_1_to_latch_low_25_port, o(24) => 
                           from_mux_2_1_to_latch_low_24_port, o(23) => 
                           from_mux_2_1_to_latch_low_23_port, o(22) => 
                           from_mux_2_1_to_latch_low_22_port, o(21) => 
                           from_mux_2_1_to_latch_low_21_port, o(20) => 
                           from_mux_2_1_to_latch_low_20_port, o(19) => 
                           from_mux_2_1_to_latch_low_19_port, o(18) => 
                           from_mux_2_1_to_latch_low_18_port, o(17) => 
                           from_mux_2_1_to_latch_low_17_port, o(16) => 
                           from_mux_2_1_to_latch_low_16_port, o(15) => 
                           from_mux_2_1_to_latch_low_15_port, o(14) => 
                           from_mux_2_1_to_latch_low_14_port, o(13) => 
                           from_mux_2_1_to_latch_low_13_port, o(12) => 
                           from_mux_2_1_to_latch_low_12_port, o(11) => 
                           from_mux_2_1_to_latch_low_11_port, o(10) => 
                           from_mux_2_1_to_latch_low_10_port, o(9) => 
                           from_mux_2_1_to_latch_low_9_port, o(8) => 
                           from_mux_2_1_to_latch_low_8_port, o(7) => 
                           from_mux_2_1_to_latch_low_7_port, o(6) => 
                           from_mux_2_1_to_latch_low_6_port, o(5) => 
                           from_mux_2_1_to_latch_low_5_port, o(4) => 
                           from_mux_2_1_to_latch_low_4_port, o(3) => 
                           from_mux_2_1_to_latch_low_3_port, o(2) => 
                           from_mux_2_1_to_latch_low_2_port, o(1) => 
                           from_mux_2_1_to_latch_low_1_port, o(0) => 
                           from_mux_2_1_to_latch_low_0_port);
   M0 : mux3_1_0 port map( operand_one(31) => operand_a(31), operand_one(30) =>
                           operand_a(30), operand_one(29) => operand_a(29), 
                           operand_one(28) => operand_a(28), operand_one(27) =>
                           operand_a(27), operand_one(26) => operand_a(26), 
                           operand_one(25) => operand_a(25), operand_one(24) =>
                           operand_a(24), operand_one(23) => operand_a(23), 
                           operand_one(22) => operand_a(22), operand_one(21) =>
                           operand_a(21), operand_one(20) => operand_a(20), 
                           operand_one(19) => operand_a(19), operand_one(18) =>
                           operand_a(18), operand_one(17) => operand_a(17), 
                           operand_one(16) => operand_a(16), operand_one(15) =>
                           operand_a(15), operand_one(14) => operand_a(14), 
                           operand_one(13) => operand_a(13), operand_one(12) =>
                           operand_a(12), operand_one(11) => operand_a(11), 
                           operand_one(10) => operand_a(10), operand_one(9) => 
                           operand_a(9), operand_one(8) => operand_a(8), 
                           operand_one(7) => operand_a(7), operand_one(6) => 
                           operand_a(6), operand_one(5) => operand_a(5), 
                           operand_one(4) => operand_a(4), operand_one(3) => 
                           operand_a(3), operand_one(2) => operand_a(2), 
                           operand_one(1) => operand_a(1), operand_one(0) => 
                           operand_a(0), operand_two(31) => forward_exe(31), 
                           operand_two(30) => forward_exe(30), operand_two(29) 
                           => forward_exe(29), operand_two(28) => 
                           forward_exe(28), operand_two(27) => forward_exe(27),
                           operand_two(26) => forward_exe(26), operand_two(25) 
                           => forward_exe(25), operand_two(24) => 
                           forward_exe(24), operand_two(23) => forward_exe(23),
                           operand_two(22) => forward_exe(22), operand_two(21) 
                           => forward_exe(21), operand_two(20) => 
                           forward_exe(20), operand_two(19) => forward_exe(19),
                           operand_two(18) => forward_exe(18), operand_two(17) 
                           => forward_exe(17), operand_two(16) => 
                           forward_exe(16), operand_two(15) => forward_exe(15),
                           operand_two(14) => forward_exe(14), operand_two(13) 
                           => forward_exe(13), operand_two(12) => 
                           forward_exe(12), operand_two(11) => forward_exe(11),
                           operand_two(10) => forward_exe(10), operand_two(9) 
                           => forward_exe(9), operand_two(8) => forward_exe(8),
                           operand_two(7) => forward_exe(7), operand_two(6) => 
                           forward_exe(6), operand_two(5) => forward_exe(5), 
                           operand_two(4) => forward_exe(4), operand_two(3) => 
                           forward_exe(3), operand_two(2) => forward_exe(2), 
                           operand_two(1) => forward_exe(1), operand_two(0) => 
                           forward_exe(0), operand_three(31) => forward_mem(31)
                           , operand_three(30) => forward_mem(30), 
                           operand_three(29) => forward_mem(29), 
                           operand_three(28) => forward_mem(28), 
                           operand_three(27) => forward_mem(27), 
                           operand_three(26) => forward_mem(26), 
                           operand_three(25) => forward_mem(25), 
                           operand_three(24) => forward_mem(24), 
                           operand_three(23) => forward_mem(23), 
                           operand_three(22) => forward_mem(22), 
                           operand_three(21) => forward_mem(21), 
                           operand_three(20) => forward_mem(20), 
                           operand_three(19) => forward_mem(19), 
                           operand_three(18) => forward_mem(18), 
                           operand_three(17) => forward_mem(17), 
                           operand_three(16) => forward_mem(16), 
                           operand_three(15) => forward_mem(15), 
                           operand_three(14) => forward_mem(14), 
                           operand_three(13) => forward_mem(13), 
                           operand_three(12) => forward_mem(12), 
                           operand_three(11) => forward_mem(11), 
                           operand_three(10) => forward_mem(10), 
                           operand_three(9) => forward_mem(9), operand_three(8)
                           => forward_mem(8), operand_three(7) => 
                           forward_mem(7), operand_three(6) => forward_mem(6), 
                           operand_three(5) => forward_mem(5), operand_three(4)
                           => forward_mem(4), operand_three(3) => 
                           forward_mem(3), operand_three(2) => forward_mem(2), 
                           operand_three(1) => forward_mem(1), operand_three(0)
                           => forward_mem(0), sel(1) => sel_mux_3_1_high_1_port
                           , sel(0) => sel_mux_3_1_high_0_port, out_res(31) => 
                           mux_to_mux_high_31_port, out_res(30) => 
                           mux_to_mux_high_30_port, out_res(29) => 
                           mux_to_mux_high_29_port, out_res(28) => 
                           mux_to_mux_high_28_port, out_res(27) => 
                           mux_to_mux_high_27_port, out_res(26) => 
                           mux_to_mux_high_26_port, out_res(25) => 
                           mux_to_mux_high_25_port, out_res(24) => 
                           mux_to_mux_high_24_port, out_res(23) => 
                           mux_to_mux_high_23_port, out_res(22) => 
                           mux_to_mux_high_22_port, out_res(21) => 
                           mux_to_mux_high_21_port, out_res(20) => 
                           mux_to_mux_high_20_port, out_res(19) => 
                           mux_to_mux_high_19_port, out_res(18) => 
                           mux_to_mux_high_18_port, out_res(17) => 
                           mux_to_mux_high_17_port, out_res(16) => 
                           mux_to_mux_high_16_port, out_res(15) => 
                           mux_to_mux_high_15_port, out_res(14) => 
                           mux_to_mux_high_14_port, out_res(13) => 
                           mux_to_mux_high_13_port, out_res(12) => 
                           mux_to_mux_high_12_port, out_res(11) => 
                           mux_to_mux_high_11_port, out_res(10) => 
                           mux_to_mux_high_10_port, out_res(9) => 
                           mux_to_mux_high_9_port, out_res(8) => 
                           mux_to_mux_high_8_port, out_res(7) => 
                           mux_to_mux_high_7_port, out_res(6) => 
                           mux_to_mux_high_6_port, out_res(5) => 
                           mux_to_mux_high_5_port, out_res(4) => 
                           mux_to_mux_high_4_port, out_res(3) => 
                           mux_to_mux_high_3_port, out_res(2) => 
                           mux_to_mux_high_2_port, out_res(1) => 
                           mux_to_mux_high_1_port, out_res(0) => 
                           mux_to_mux_high_0_port);
   M1 : mux3_1_1 port map( operand_one(31) => operand_b(31), operand_one(30) =>
                           operand_b(30), operand_one(29) => operand_b(29), 
                           operand_one(28) => operand_b(28), operand_one(27) =>
                           operand_b(27), operand_one(26) => operand_b(26), 
                           operand_one(25) => operand_b(25), operand_one(24) =>
                           operand_b(24), operand_one(23) => operand_b(23), 
                           operand_one(22) => operand_b(22), operand_one(21) =>
                           operand_b(21), operand_one(20) => operand_b(20), 
                           operand_one(19) => operand_b(19), operand_one(18) =>
                           operand_b(18), operand_one(17) => operand_b(17), 
                           operand_one(16) => operand_b(16), operand_one(15) =>
                           operand_b(15), operand_one(14) => operand_b(14), 
                           operand_one(13) => operand_b(13), operand_one(12) =>
                           operand_b(12), operand_one(11) => operand_b(11), 
                           operand_one(10) => operand_b(10), operand_one(9) => 
                           operand_b(9), operand_one(8) => operand_b(8), 
                           operand_one(7) => operand_b(7), operand_one(6) => 
                           operand_b(6), operand_one(5) => operand_b(5), 
                           operand_one(4) => operand_b(4), operand_one(3) => 
                           operand_b(3), operand_one(2) => operand_b(2), 
                           operand_one(1) => operand_b(1), operand_one(0) => 
                           operand_b(0), operand_two(31) => forward_exe(31), 
                           operand_two(30) => forward_exe(30), operand_two(29) 
                           => forward_exe(29), operand_two(28) => 
                           forward_exe(28), operand_two(27) => forward_exe(27),
                           operand_two(26) => forward_exe(26), operand_two(25) 
                           => forward_exe(25), operand_two(24) => 
                           forward_exe(24), operand_two(23) => forward_exe(23),
                           operand_two(22) => forward_exe(22), operand_two(21) 
                           => forward_exe(21), operand_two(20) => 
                           forward_exe(20), operand_two(19) => forward_exe(19),
                           operand_two(18) => forward_exe(18), operand_two(17) 
                           => forward_exe(17), operand_two(16) => 
                           forward_exe(16), operand_two(15) => forward_exe(15),
                           operand_two(14) => forward_exe(14), operand_two(13) 
                           => forward_exe(13), operand_two(12) => 
                           forward_exe(12), operand_two(11) => forward_exe(11),
                           operand_two(10) => forward_exe(10), operand_two(9) 
                           => forward_exe(9), operand_two(8) => forward_exe(8),
                           operand_two(7) => forward_exe(7), operand_two(6) => 
                           forward_exe(6), operand_two(5) => forward_exe(5), 
                           operand_two(4) => forward_exe(4), operand_two(3) => 
                           forward_exe(3), operand_two(2) => forward_exe(2), 
                           operand_two(1) => forward_exe(1), operand_two(0) => 
                           forward_exe(0), operand_three(31) => forward_mem(31)
                           , operand_three(30) => forward_mem(30), 
                           operand_three(29) => forward_mem(29), 
                           operand_three(28) => forward_mem(28), 
                           operand_three(27) => forward_mem(27), 
                           operand_three(26) => forward_mem(26), 
                           operand_three(25) => forward_mem(25), 
                           operand_three(24) => forward_mem(24), 
                           operand_three(23) => forward_mem(23), 
                           operand_three(22) => forward_mem(22), 
                           operand_three(21) => forward_mem(21), 
                           operand_three(20) => forward_mem(20), 
                           operand_three(19) => forward_mem(19), 
                           operand_three(18) => forward_mem(18), 
                           operand_three(17) => forward_mem(17), 
                           operand_three(16) => forward_mem(16), 
                           operand_three(15) => forward_mem(15), 
                           operand_three(14) => forward_mem(14), 
                           operand_three(13) => forward_mem(13), 
                           operand_three(12) => forward_mem(12), 
                           operand_three(11) => forward_mem(11), 
                           operand_three(10) => forward_mem(10), 
                           operand_three(9) => forward_mem(9), operand_three(8)
                           => forward_mem(8), operand_three(7) => 
                           forward_mem(7), operand_three(6) => forward_mem(6), 
                           operand_three(5) => forward_mem(5), operand_three(4)
                           => forward_mem(4), operand_three(3) => 
                           forward_mem(3), operand_three(2) => forward_mem(2), 
                           operand_three(1) => forward_mem(1), operand_three(0)
                           => forward_mem(0), sel(1) => sel_mux_3_1_low_1_port,
                           sel(0) => sel_mux_3_1_low_0_port, out_res(31) => 
                           mux_to_mux_low_31_port, out_res(30) => 
                           mux_to_mux_low_30_port, out_res(29) => 
                           mux_to_mux_low_29_port, out_res(28) => 
                           mux_to_mux_low_28_port, out_res(27) => 
                           mux_to_mux_low_27_port, out_res(26) => 
                           mux_to_mux_low_26_port, out_res(25) => 
                           mux_to_mux_low_25_port, out_res(24) => 
                           mux_to_mux_low_24_port, out_res(23) => 
                           mux_to_mux_low_23_port, out_res(22) => 
                           mux_to_mux_low_22_port, out_res(21) => 
                           mux_to_mux_low_21_port, out_res(20) => 
                           mux_to_mux_low_20_port, out_res(19) => 
                           mux_to_mux_low_19_port, out_res(18) => 
                           mux_to_mux_low_18_port, out_res(17) => 
                           mux_to_mux_low_17_port, out_res(16) => 
                           mux_to_mux_low_16_port, out_res(15) => 
                           mux_to_mux_low_15_port, out_res(14) => 
                           mux_to_mux_low_14_port, out_res(13) => 
                           mux_to_mux_low_13_port, out_res(12) => 
                           mux_to_mux_low_12_port, out_res(11) => 
                           mux_to_mux_low_11_port, out_res(10) => 
                           mux_to_mux_low_10_port, out_res(9) => 
                           mux_to_mux_low_9_port, out_res(8) => 
                           mux_to_mux_low_8_port, out_res(7) => 
                           mux_to_mux_low_7_port, out_res(6) => 
                           mux_to_mux_low_6_port, out_res(5) => 
                           mux_to_mux_low_5_port, out_res(4) => 
                           mux_to_mux_low_4_port, out_res(3) => 
                           mux_to_mux_low_3_port, out_res(2) => 
                           mux_to_mux_low_2_port, out_res(1) => 
                           mux_to_mux_low_1_port, out_res(0) => 
                           mux_to_mux_low_0_port);
   n4 <= '0';

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity memoryUnit is

   port( clock, reset, enable : in std_logic;  alu_result, data_from_memory : 
         in std_logic_vector (31 downto 0);  EX_MEM_Rd : in std_logic_vector (4
         downto 0);  address_memory, data_op1, data_op2 : out std_logic_vector 
         (31 downto 0);  MEM_WB_Rd : out std_logic_vector (4 downto 0));

end memoryUnit;

architecture SYN_Behavioral of memoryUnit is

   component regWithEnable_7
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component regWithEnable_8
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component regWithEnable_5bit_0
      port( input : in std_logic_vector (4 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (4 downto 0));
   end component;

begin
   address_memory <= ( alu_result(31), alu_result(30), alu_result(29), 
      alu_result(28), alu_result(27), alu_result(26), alu_result(25), 
      alu_result(24), alu_result(23), alu_result(22), alu_result(21), 
      alu_result(20), alu_result(19), alu_result(18), alu_result(17), 
      alu_result(16), alu_result(15), alu_result(14), alu_result(13), 
      alu_result(12), alu_result(11), alu_result(10), alu_result(9), 
      alu_result(8), alu_result(7), alu_result(6), alu_result(5), alu_result(4)
      , alu_result(3), alu_result(2), alu_result(1), alu_result(0) );
   
   RE : regWithEnable_5bit_0 port map( input(4) => EX_MEM_Rd(4), input(3) => 
                           EX_MEM_Rd(3), input(2) => EX_MEM_Rd(2), input(1) => 
                           EX_MEM_Rd(1), input(0) => EX_MEM_Rd(0), en => enable
                           , clock => clock, reset => reset, output(4) => 
                           MEM_WB_Rd(4), output(3) => MEM_WB_Rd(3), output(2) 
                           => MEM_WB_Rd(2), output(1) => MEM_WB_Rd(1), 
                           output(0) => MEM_WB_Rd(0));
   RE_1 : regWithEnable_8 port map( input(31) => data_from_memory(31), 
                           input(30) => data_from_memory(30), input(29) => 
                           data_from_memory(29), input(28) => 
                           data_from_memory(28), input(27) => 
                           data_from_memory(27), input(26) => 
                           data_from_memory(26), input(25) => 
                           data_from_memory(25), input(24) => 
                           data_from_memory(24), input(23) => 
                           data_from_memory(23), input(22) => 
                           data_from_memory(22), input(21) => 
                           data_from_memory(21), input(20) => 
                           data_from_memory(20), input(19) => 
                           data_from_memory(19), input(18) => 
                           data_from_memory(18), input(17) => 
                           data_from_memory(17), input(16) => 
                           data_from_memory(16), input(15) => 
                           data_from_memory(15), input(14) => 
                           data_from_memory(14), input(13) => 
                           data_from_memory(13), input(12) => 
                           data_from_memory(12), input(11) => 
                           data_from_memory(11), input(10) => 
                           data_from_memory(10), input(9) => 
                           data_from_memory(9), input(8) => data_from_memory(8)
                           , input(7) => data_from_memory(7), input(6) => 
                           data_from_memory(6), input(5) => data_from_memory(5)
                           , input(4) => data_from_memory(4), input(3) => 
                           data_from_memory(3), input(2) => data_from_memory(2)
                           , input(1) => data_from_memory(1), input(0) => 
                           data_from_memory(0), en => enable, clock => clock, 
                           reset => reset, output(31) => data_op1(31), 
                           output(30) => data_op1(30), output(29) => 
                           data_op1(29), output(28) => data_op1(28), output(27)
                           => data_op1(27), output(26) => data_op1(26), 
                           output(25) => data_op1(25), output(24) => 
                           data_op1(24), output(23) => data_op1(23), output(22)
                           => data_op1(22), output(21) => data_op1(21), 
                           output(20) => data_op1(20), output(19) => 
                           data_op1(19), output(18) => data_op1(18), output(17)
                           => data_op1(17), output(16) => data_op1(16), 
                           output(15) => data_op1(15), output(14) => 
                           data_op1(14), output(13) => data_op1(13), output(12)
                           => data_op1(12), output(11) => data_op1(11), 
                           output(10) => data_op1(10), output(9) => data_op1(9)
                           , output(8) => data_op1(8), output(7) => data_op1(7)
                           , output(6) => data_op1(6), output(5) => data_op1(5)
                           , output(4) => data_op1(4), output(3) => data_op1(3)
                           , output(2) => data_op1(2), output(1) => data_op1(1)
                           , output(0) => data_op1(0));
   RE_2 : regWithEnable_7 port map( input(31) => alu_result(31), input(30) => 
                           alu_result(30), input(29) => alu_result(29), 
                           input(28) => alu_result(28), input(27) => 
                           alu_result(27), input(26) => alu_result(26), 
                           input(25) => alu_result(25), input(24) => 
                           alu_result(24), input(23) => alu_result(23), 
                           input(22) => alu_result(22), input(21) => 
                           alu_result(21), input(20) => alu_result(20), 
                           input(19) => alu_result(19), input(18) => 
                           alu_result(18), input(17) => alu_result(17), 
                           input(16) => alu_result(16), input(15) => 
                           alu_result(15), input(14) => alu_result(14), 
                           input(13) => alu_result(13), input(12) => 
                           alu_result(12), input(11) => alu_result(11), 
                           input(10) => alu_result(10), input(9) => 
                           alu_result(9), input(8) => alu_result(8), input(7) 
                           => alu_result(7), input(6) => alu_result(6), 
                           input(5) => alu_result(5), input(4) => alu_result(4)
                           , input(3) => alu_result(3), input(2) => 
                           alu_result(2), input(1) => alu_result(1), input(0) 
                           => alu_result(0), en => enable, clock => clock, 
                           reset => reset, output(31) => data_op2(31), 
                           output(30) => data_op2(30), output(29) => 
                           data_op2(29), output(28) => data_op2(28), output(27)
                           => data_op2(27), output(26) => data_op2(26), 
                           output(25) => data_op2(25), output(24) => 
                           data_op2(24), output(23) => data_op2(23), output(22)
                           => data_op2(22), output(21) => data_op2(21), 
                           output(20) => data_op2(20), output(19) => 
                           data_op2(19), output(18) => data_op2(18), output(17)
                           => data_op2(17), output(16) => data_op2(16), 
                           output(15) => data_op2(15), output(14) => 
                           data_op2(14), output(13) => data_op2(13), output(12)
                           => data_op2(12), output(11) => data_op2(11), 
                           output(10) => data_op2(10), output(9) => data_op2(9)
                           , output(8) => data_op2(8), output(7) => data_op2(7)
                           , output(6) => data_op2(6), output(5) => data_op2(5)
                           , output(4) => data_op2(4), output(3) => data_op2(3)
                           , output(2) => data_op2(2), output(1) => data_op2(1)
                           , output(0) => data_op2(0));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity writeBacKUnit is

   port( clock, reset, enable, sel_4 : in std_logic;  data_from_memory, 
         data_from_alu : in std_logic_vector (31 downto 0);  write_back_value, 
         debug : out std_logic_vector (31 downto 0));

end writeBacKUnit;

architecture SYN_Behavioral of writeBacKUnit is

   component regWithEnable_0
      port( input : in std_logic_vector (31 downto 0);  en, clock, reset : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux2X1_0
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  o :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal write_back_value_31_port, write_back_value_30_port, 
      write_back_value_29_port, write_back_value_28_port, 
      write_back_value_27_port, write_back_value_26_port, 
      write_back_value_25_port, write_back_value_24_port, 
      write_back_value_23_port, write_back_value_22_port, 
      write_back_value_21_port, write_back_value_20_port, 
      write_back_value_19_port, write_back_value_18_port, 
      write_back_value_17_port, write_back_value_16_port, 
      write_back_value_15_port, write_back_value_14_port, 
      write_back_value_13_port, write_back_value_12_port, 
      write_back_value_11_port, write_back_value_10_port, 
      write_back_value_9_port, write_back_value_8_port, write_back_value_7_port
      , write_back_value_6_port, write_back_value_5_port, 
      write_back_value_4_port, write_back_value_3_port, write_back_value_2_port
      , write_back_value_1_port, write_back_value_0_port : std_logic;

begin
   write_back_value <= ( write_back_value_31_port, write_back_value_30_port, 
      write_back_value_29_port, write_back_value_28_port, 
      write_back_value_27_port, write_back_value_26_port, 
      write_back_value_25_port, write_back_value_24_port, 
      write_back_value_23_port, write_back_value_22_port, 
      write_back_value_21_port, write_back_value_20_port, 
      write_back_value_19_port, write_back_value_18_port, 
      write_back_value_17_port, write_back_value_16_port, 
      write_back_value_15_port, write_back_value_14_port, 
      write_back_value_13_port, write_back_value_12_port, 
      write_back_value_11_port, write_back_value_10_port, 
      write_back_value_9_port, write_back_value_8_port, write_back_value_7_port
      , write_back_value_6_port, write_back_value_5_port, 
      write_back_value_4_port, write_back_value_3_port, write_back_value_2_port
      , write_back_value_1_port, write_back_value_0_port );
   
   M0 : Mux2X1_0 port map( a(31) => data_from_memory(31), a(30) => 
                           data_from_memory(30), a(29) => data_from_memory(29),
                           a(28) => data_from_memory(28), a(27) => 
                           data_from_memory(27), a(26) => data_from_memory(26),
                           a(25) => data_from_memory(25), a(24) => 
                           data_from_memory(24), a(23) => data_from_memory(23),
                           a(22) => data_from_memory(22), a(21) => 
                           data_from_memory(21), a(20) => data_from_memory(20),
                           a(19) => data_from_memory(19), a(18) => 
                           data_from_memory(18), a(17) => data_from_memory(17),
                           a(16) => data_from_memory(16), a(15) => 
                           data_from_memory(15), a(14) => data_from_memory(14),
                           a(13) => data_from_memory(13), a(12) => 
                           data_from_memory(12), a(11) => data_from_memory(11),
                           a(10) => data_from_memory(10), a(9) => 
                           data_from_memory(9), a(8) => data_from_memory(8), 
                           a(7) => data_from_memory(7), a(6) => 
                           data_from_memory(6), a(5) => data_from_memory(5), 
                           a(4) => data_from_memory(4), a(3) => 
                           data_from_memory(3), a(2) => data_from_memory(2), 
                           a(1) => data_from_memory(1), a(0) => 
                           data_from_memory(0), b(31) => data_from_alu(31), 
                           b(30) => data_from_alu(30), b(29) => 
                           data_from_alu(29), b(28) => data_from_alu(28), b(27)
                           => data_from_alu(27), b(26) => data_from_alu(26), 
                           b(25) => data_from_alu(25), b(24) => 
                           data_from_alu(24), b(23) => data_from_alu(23), b(22)
                           => data_from_alu(22), b(21) => data_from_alu(21), 
                           b(20) => data_from_alu(20), b(19) => 
                           data_from_alu(19), b(18) => data_from_alu(18), b(17)
                           => data_from_alu(17), b(16) => data_from_alu(16), 
                           b(15) => data_from_alu(15), b(14) => 
                           data_from_alu(14), b(13) => data_from_alu(13), b(12)
                           => data_from_alu(12), b(11) => data_from_alu(11), 
                           b(10) => data_from_alu(10), b(9) => data_from_alu(9)
                           , b(8) => data_from_alu(8), b(7) => data_from_alu(7)
                           , b(6) => data_from_alu(6), b(5) => data_from_alu(5)
                           , b(4) => data_from_alu(4), b(3) => data_from_alu(3)
                           , b(2) => data_from_alu(2), b(1) => data_from_alu(1)
                           , b(0) => data_from_alu(0), sel => sel_4, o(31) => 
                           write_back_value_31_port, o(30) => 
                           write_back_value_30_port, o(29) => 
                           write_back_value_29_port, o(28) => 
                           write_back_value_28_port, o(27) => 
                           write_back_value_27_port, o(26) => 
                           write_back_value_26_port, o(25) => 
                           write_back_value_25_port, o(24) => 
                           write_back_value_24_port, o(23) => 
                           write_back_value_23_port, o(22) => 
                           write_back_value_22_port, o(21) => 
                           write_back_value_21_port, o(20) => 
                           write_back_value_20_port, o(19) => 
                           write_back_value_19_port, o(18) => 
                           write_back_value_18_port, o(17) => 
                           write_back_value_17_port, o(16) => 
                           write_back_value_16_port, o(15) => 
                           write_back_value_15_port, o(14) => 
                           write_back_value_14_port, o(13) => 
                           write_back_value_13_port, o(12) => 
                           write_back_value_12_port, o(11) => 
                           write_back_value_11_port, o(10) => 
                           write_back_value_10_port, o(9) => 
                           write_back_value_9_port, o(8) => 
                           write_back_value_8_port, o(7) => 
                           write_back_value_7_port, o(6) => 
                           write_back_value_6_port, o(5) => 
                           write_back_value_5_port, o(4) => 
                           write_back_value_4_port, o(3) => 
                           write_back_value_3_port, o(2) => 
                           write_back_value_2_port, o(1) => 
                           write_back_value_1_port, o(0) => 
                           write_back_value_0_port);
   RE_DEBUG : regWithEnable_0 port map( input(31) => write_back_value_31_port, 
                           input(30) => write_back_value_30_port, input(29) => 
                           write_back_value_29_port, input(28) => 
                           write_back_value_28_port, input(27) => 
                           write_back_value_27_port, input(26) => 
                           write_back_value_26_port, input(25) => 
                           write_back_value_25_port, input(24) => 
                           write_back_value_24_port, input(23) => 
                           write_back_value_23_port, input(22) => 
                           write_back_value_22_port, input(21) => 
                           write_back_value_21_port, input(20) => 
                           write_back_value_20_port, input(19) => 
                           write_back_value_19_port, input(18) => 
                           write_back_value_18_port, input(17) => 
                           write_back_value_17_port, input(16) => 
                           write_back_value_16_port, input(15) => 
                           write_back_value_15_port, input(14) => 
                           write_back_value_14_port, input(13) => 
                           write_back_value_13_port, input(12) => 
                           write_back_value_12_port, input(11) => 
                           write_back_value_11_port, input(10) => 
                           write_back_value_10_port, input(9) => 
                           write_back_value_9_port, input(8) => 
                           write_back_value_8_port, input(7) => 
                           write_back_value_7_port, input(6) => 
                           write_back_value_6_port, input(5) => 
                           write_back_value_5_port, input(4) => 
                           write_back_value_4_port, input(3) => 
                           write_back_value_3_port, input(2) => 
                           write_back_value_2_port, input(1) => 
                           write_back_value_1_port, input(0) => 
                           write_back_value_0_port, en => enable, clock => 
                           clock, reset => reset, output(31) => debug(31), 
                           output(30) => debug(30), output(29) => debug(29), 
                           output(28) => debug(28), output(27) => debug(27), 
                           output(26) => debug(26), output(25) => debug(25), 
                           output(24) => debug(24), output(23) => debug(23), 
                           output(22) => debug(22), output(21) => debug(21), 
                           output(20) => debug(20), output(19) => debug(19), 
                           output(18) => debug(18), output(17) => debug(17), 
                           output(16) => debug(16), output(15) => debug(15), 
                           output(14) => debug(14), output(13) => debug(13), 
                           output(12) => debug(12), output(11) => debug(11), 
                           output(10) => debug(10), output(9) => debug(9), 
                           output(8) => debug(8), output(7) => debug(7), 
                           output(6) => debug(6), output(5) => debug(5), 
                           output(4) => debug(4), output(3) => debug(3), 
                           output(2) => debug(2), output(1) => debug(1), 
                           output(0) => debug(0));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_dataPath.all;

entity dataPath is

   port( sel0, sel1, sel2, sel3, sel4, sel_ext, en1, en2, en3, en4, en5, en6, 
         en7, clock, reset, hazard_condition : in std_logic;  func : in 
         std_logic_vector (10 downto 0);  EX_MEM_write, MEM_WB_write : in 
         std_logic;  from_instruction_memory, datain : in std_logic_vector (31 
         downto 0);  hazard_detected, jump : out std_logic;  pc_to_im, 
         instruction, address_data_memory, dataout, debug : out 
         std_logic_vector (31 downto 0));

end dataPath;

architecture SYN_Structural of dataPath is

   component fetchUnit
      port( sel0, en0, clock, reset : in std_logic;  fromInstructionMemory, 
            next_PC : in std_logic_vector (31 downto 0);  PcToInstructionMemory
            , InstructionToDecode, pcToDecode : out std_logic_vector (31 downto
            0));
   end component;
   
   component decodeUnit
      port( clock, reset, en1, read_enable_portA, read_enable_portB, 
            write_enable_portW : in std_logic;  instructionWord : in 
            std_logic_vector (31 downto 0);  ID_EX_MemRead : in std_logic;  
            ID_EX_RT_Address : in std_logic_vector (4 downto 0);  writeData : 
            in std_logic_vector (31 downto 0);  writeAddress : in 
            std_logic_vector (4 downto 0);  pc : in std_logic_vector (31 downto
            0);  sel_ext, multi_cycle_operation : in std_logic;  
            enable_signal_PC_IF_ID, selectNop : out std_logic;  outRT, outRD, 
            outRS : out std_logic_vector (4 downto 0);  outIMM, outPC, outA, 
            outB : out std_logic_vector (31 downto 0));
   end component;
   
   component executionUnit
      port( clock, reset : in std_logic;  operand_a, operand_b, operand_imm, 
            operand_pc, forward_exe, forward_mem : in std_logic_vector (31 
            downto 0);  EX_MEM_write, MEM_WB_write : in std_logic;  MEM_WB_rd, 
            ID_EX_Rd, ID_EX_Rs, ID_EX_Rt : in std_logic_vector (4 downto 0);  
            enable, sel_1, sel_2, sel_3 : in std_logic;  func : in 
            std_logic_vector (10 downto 0);  EX_MEM_rd : inout std_logic_vector
            (4 downto 0);  out_res_operand_one, out_res_operand_two, next_pc : 
            out std_logic_vector (31 downto 0);  jump, multi_cycle_operation : 
            out std_logic);
   end component;
   
   component memoryUnit
      port( clock, reset, enable : in std_logic;  alu_result, data_from_memory 
            : in std_logic_vector (31 downto 0);  EX_MEM_Rd : in 
            std_logic_vector (4 downto 0);  address_memory, data_op1, data_op2 
            : out std_logic_vector (31 downto 0);  MEM_WB_Rd : out 
            std_logic_vector (4 downto 0));
   end component;
   
   component writeBacKUnit
      port( clock, reset, enable, sel_4 : in std_logic;  data_from_memory, 
            data_from_alu : in std_logic_vector (31 downto 0);  
            write_back_value, debug : out std_logic_vector (31 downto 0));
   end component;
   
   signal instruction_31_port, instruction_30_port, instruction_29_port, 
      instruction_28_port, instruction_27_port, instruction_26_port, 
      instruction_25_port, instruction_24_port, instruction_23_port, 
      instruction_22_port, instruction_21_port, instruction_20_port, 
      instruction_19_port, instruction_18_port, instruction_17_port, 
      instruction_16_port, instruction_15_port, instruction_14_port, 
      instruction_13_port, instruction_12_port, instruction_11_port, 
      instruction_10_port, instruction_9_port, instruction_8_port, 
      instruction_7_port, instruction_6_port, instruction_5_port, 
      instruction_4_port, instruction_3_port, instruction_2_port, 
      instruction_1_port, instruction_0_port, write_back_op1_31_port, 
      write_back_op1_30_port, write_back_op1_29_port, write_back_op1_28_port, 
      write_back_op1_27_port, write_back_op1_26_port, write_back_op1_25_port, 
      write_back_op1_24_port, write_back_op1_23_port, write_back_op1_22_port, 
      write_back_op1_21_port, write_back_op1_20_port, write_back_op1_19_port, 
      write_back_op1_18_port, write_back_op1_17_port, write_back_op1_16_port, 
      write_back_op1_15_port, write_back_op1_14_port, write_back_op1_13_port, 
      write_back_op1_12_port, write_back_op1_11_port, write_back_op1_10_port, 
      write_back_op1_9_port, write_back_op1_8_port, write_back_op1_7_port, 
      write_back_op1_6_port, write_back_op1_5_port, write_back_op1_4_port, 
      write_back_op1_3_port, write_back_op1_2_port, write_back_op1_1_port, 
      write_back_op1_0_port, write_back_op2_31_port, write_back_op2_30_port, 
      write_back_op2_29_port, write_back_op2_28_port, write_back_op2_27_port, 
      write_back_op2_26_port, write_back_op2_25_port, write_back_op2_24_port, 
      write_back_op2_23_port, write_back_op2_22_port, write_back_op2_21_port, 
      write_back_op2_20_port, write_back_op2_19_port, write_back_op2_18_port, 
      write_back_op2_17_port, write_back_op2_16_port, write_back_op2_15_port, 
      write_back_op2_14_port, write_back_op2_13_port, write_back_op2_12_port, 
      write_back_op2_11_port, write_back_op2_10_port, write_back_op2_9_port, 
      write_back_op2_8_port, write_back_op2_7_port, write_back_op2_6_port, 
      write_back_op2_5_port, write_back_op2_4_port, write_back_op2_3_port, 
      write_back_op2_2_port, write_back_op2_1_port, write_back_op2_0_port, 
      forward_mem_31_port, forward_mem_30_port, forward_mem_29_port, 
      forward_mem_28_port, forward_mem_27_port, forward_mem_26_port, 
      forward_mem_25_port, forward_mem_24_port, forward_mem_23_port, 
      forward_mem_22_port, forward_mem_21_port, forward_mem_20_port, 
      forward_mem_19_port, forward_mem_18_port, forward_mem_17_port, 
      forward_mem_16_port, forward_mem_15_port, forward_mem_14_port, 
      forward_mem_13_port, forward_mem_12_port, forward_mem_11_port, 
      forward_mem_10_port, forward_mem_9_port, forward_mem_8_port, 
      forward_mem_7_port, forward_mem_6_port, forward_mem_5_port, 
      forward_mem_4_port, forward_mem_3_port, forward_mem_2_port, 
      forward_mem_1_port, forward_mem_0_port, operand_res_alu_31_port, 
      operand_res_alu_30_port, operand_res_alu_29_port, operand_res_alu_28_port
      , operand_res_alu_27_port, operand_res_alu_26_port, 
      operand_res_alu_25_port, operand_res_alu_24_port, operand_res_alu_23_port
      , operand_res_alu_22_port, operand_res_alu_21_port, 
      operand_res_alu_20_port, operand_res_alu_19_port, operand_res_alu_18_port
      , operand_res_alu_17_port, operand_res_alu_16_port, 
      operand_res_alu_15_port, operand_res_alu_14_port, operand_res_alu_13_port
      , operand_res_alu_12_port, operand_res_alu_11_port, 
      operand_res_alu_10_port, operand_res_alu_9_port, operand_res_alu_8_port, 
      operand_res_alu_7_port, operand_res_alu_6_port, operand_res_alu_5_port, 
      operand_res_alu_4_port, operand_res_alu_3_port, operand_res_alu_2_port, 
      operand_res_alu_1_port, operand_res_alu_0_port, EX_MEM_RD_4_port, 
      EX_MEM_RD_3_port, EX_MEM_RD_2_port, EX_MEM_RD_1_port, EX_MEM_RD_0_port, 
      MEM_WB_RD_4_port, MEM_WB_RD_3_port, MEM_WB_RD_2_port, MEM_WB_RD_1_port, 
      MEM_WB_RD_0_port, operand_A_31_port, operand_A_30_port, operand_A_29_port
      , operand_A_28_port, operand_A_27_port, operand_A_26_port, 
      operand_A_25_port, operand_A_24_port, operand_A_23_port, 
      operand_A_22_port, operand_A_21_port, operand_A_20_port, 
      operand_A_19_port, operand_A_18_port, operand_A_17_port, 
      operand_A_16_port, operand_A_15_port, operand_A_14_port, 
      operand_A_13_port, operand_A_12_port, operand_A_11_port, 
      operand_A_10_port, operand_A_9_port, operand_A_8_port, operand_A_7_port, 
      operand_A_6_port, operand_A_5_port, operand_A_4_port, operand_A_3_port, 
      operand_A_2_port, operand_A_1_port, operand_A_0_port, operand_B_31_port, 
      operand_B_30_port, operand_B_29_port, operand_B_28_port, 
      operand_B_27_port, operand_B_26_port, operand_B_25_port, 
      operand_B_24_port, operand_B_23_port, operand_B_22_port, 
      operand_B_21_port, operand_B_20_port, operand_B_19_port, 
      operand_B_18_port, operand_B_17_port, operand_B_16_port, 
      operand_B_15_port, operand_B_14_port, operand_B_13_port, 
      operand_B_12_port, operand_B_11_port, operand_B_10_port, operand_B_9_port
      , operand_B_8_port, operand_B_7_port, operand_B_6_port, operand_B_5_port,
      operand_B_4_port, operand_B_3_port, operand_B_2_port, operand_B_1_port, 
      operand_B_0_port, operand_IMM_31_port, operand_IMM_30_port, 
      operand_IMM_29_port, operand_IMM_28_port, operand_IMM_27_port, 
      operand_IMM_26_port, operand_IMM_25_port, operand_IMM_24_port, 
      operand_IMM_23_port, operand_IMM_22_port, operand_IMM_21_port, 
      operand_IMM_20_port, operand_IMM_19_port, operand_IMM_18_port, 
      operand_IMM_17_port, operand_IMM_16_port, operand_IMM_15_port, 
      operand_IMM_14_port, operand_IMM_13_port, operand_IMM_12_port, 
      operand_IMM_11_port, operand_IMM_10_port, operand_IMM_9_port, 
      operand_IMM_8_port, operand_IMM_7_port, operand_IMM_6_port, 
      operand_IMM_5_port, operand_IMM_4_port, operand_IMM_3_port, 
      operand_IMM_2_port, operand_IMM_1_port, operand_IMM_0_port, 
      operand_PC_31_port, operand_PC_30_port, operand_PC_29_port, 
      operand_PC_28_port, operand_PC_27_port, operand_PC_26_port, 
      operand_PC_25_port, operand_PC_24_port, operand_PC_23_port, 
      operand_PC_22_port, operand_PC_21_port, operand_PC_20_port, 
      operand_PC_19_port, operand_PC_18_port, operand_PC_17_port, 
      operand_PC_16_port, operand_PC_15_port, operand_PC_14_port, 
      operand_PC_13_port, operand_PC_12_port, operand_PC_11_port, 
      operand_PC_10_port, operand_PC_9_port, operand_PC_8_port, 
      operand_PC_7_port, operand_PC_6_port, operand_PC_5_port, 
      operand_PC_4_port, operand_PC_3_port, operand_PC_2_port, 
      operand_PC_1_port, operand_PC_0_port, ID_EX_Rd_4_port, ID_EX_Rd_3_port, 
      ID_EX_Rd_2_port, ID_EX_Rd_1_port, ID_EX_Rd_0_port, ID_EX_Rs_4_port, 
      ID_EX_Rs_3_port, ID_EX_Rs_2_port, ID_EX_Rs_1_port, ID_EX_Rs_0_port, 
      ID_EX_Rt_4_port, ID_EX_Rt_3_port, ID_EX_Rt_2_port, ID_EX_Rt_1_port, 
      ID_EX_Rt_0_port, next_pc_31_port, next_pc_30_port, next_pc_29_port, 
      next_pc_28_port, next_pc_27_port, next_pc_26_port, next_pc_25_port, 
      next_pc_24_port, next_pc_23_port, next_pc_22_port, next_pc_21_port, 
      next_pc_20_port, next_pc_19_port, next_pc_18_port, next_pc_17_port, 
      next_pc_16_port, next_pc_15_port, next_pc_14_port, next_pc_13_port, 
      next_pc_12_port, next_pc_11_port, next_pc_10_port, next_pc_9_port, 
      next_pc_8_port, next_pc_7_port, next_pc_6_port, next_pc_5_port, 
      next_pc_4_port, next_pc_3_port, next_pc_2_port, next_pc_1_port, 
      next_pc_0_port, multi_cycle_operation, NPC_to_decode_31_port, 
      NPC_to_decode_30_port, NPC_to_decode_29_port, NPC_to_decode_28_port, 
      NPC_to_decode_27_port, NPC_to_decode_26_port, NPC_to_decode_25_port, 
      NPC_to_decode_24_port, NPC_to_decode_23_port, NPC_to_decode_22_port, 
      NPC_to_decode_21_port, NPC_to_decode_20_port, NPC_to_decode_19_port, 
      NPC_to_decode_18_port, NPC_to_decode_17_port, NPC_to_decode_16_port, 
      NPC_to_decode_15_port, NPC_to_decode_14_port, NPC_to_decode_13_port, 
      NPC_to_decode_12_port, NPC_to_decode_11_port, NPC_to_decode_10_port, 
      NPC_to_decode_9_port, NPC_to_decode_8_port, NPC_to_decode_7_port, 
      NPC_to_decode_6_port, NPC_to_decode_5_port, NPC_to_decode_4_port, 
      NPC_to_decode_3_port, NPC_to_decode_2_port, NPC_to_decode_1_port, 
      NPC_to_decode_0_port, disable_fetch_register : std_logic;

begin
   instruction <= ( instruction_31_port, instruction_30_port, 
      instruction_29_port, instruction_28_port, instruction_27_port, 
      instruction_26_port, instruction_25_port, instruction_24_port, 
      instruction_23_port, instruction_22_port, instruction_21_port, 
      instruction_20_port, instruction_19_port, instruction_18_port, 
      instruction_17_port, instruction_16_port, instruction_15_port, 
      instruction_14_port, instruction_13_port, instruction_12_port, 
      instruction_11_port, instruction_10_port, instruction_9_port, 
      instruction_8_port, instruction_7_port, instruction_6_port, 
      instruction_5_port, instruction_4_port, instruction_3_port, 
      instruction_2_port, instruction_1_port, instruction_0_port );
   
   WB : writeBacKUnit port map( clock => clock, reset => reset, enable => en7, 
                           sel_4 => sel4, data_from_memory(31) => 
                           write_back_op1_31_port, data_from_memory(30) => 
                           write_back_op1_30_port, data_from_memory(29) => 
                           write_back_op1_29_port, data_from_memory(28) => 
                           write_back_op1_28_port, data_from_memory(27) => 
                           write_back_op1_27_port, data_from_memory(26) => 
                           write_back_op1_26_port, data_from_memory(25) => 
                           write_back_op1_25_port, data_from_memory(24) => 
                           write_back_op1_24_port, data_from_memory(23) => 
                           write_back_op1_23_port, data_from_memory(22) => 
                           write_back_op1_22_port, data_from_memory(21) => 
                           write_back_op1_21_port, data_from_memory(20) => 
                           write_back_op1_20_port, data_from_memory(19) => 
                           write_back_op1_19_port, data_from_memory(18) => 
                           write_back_op1_18_port, data_from_memory(17) => 
                           write_back_op1_17_port, data_from_memory(16) => 
                           write_back_op1_16_port, data_from_memory(15) => 
                           write_back_op1_15_port, data_from_memory(14) => 
                           write_back_op1_14_port, data_from_memory(13) => 
                           write_back_op1_13_port, data_from_memory(12) => 
                           write_back_op1_12_port, data_from_memory(11) => 
                           write_back_op1_11_port, data_from_memory(10) => 
                           write_back_op1_10_port, data_from_memory(9) => 
                           write_back_op1_9_port, data_from_memory(8) => 
                           write_back_op1_8_port, data_from_memory(7) => 
                           write_back_op1_7_port, data_from_memory(6) => 
                           write_back_op1_6_port, data_from_memory(5) => 
                           write_back_op1_5_port, data_from_memory(4) => 
                           write_back_op1_4_port, data_from_memory(3) => 
                           write_back_op1_3_port, data_from_memory(2) => 
                           write_back_op1_2_port, data_from_memory(1) => 
                           write_back_op1_1_port, data_from_memory(0) => 
                           write_back_op1_0_port, data_from_alu(31) => 
                           write_back_op2_31_port, data_from_alu(30) => 
                           write_back_op2_30_port, data_from_alu(29) => 
                           write_back_op2_29_port, data_from_alu(28) => 
                           write_back_op2_28_port, data_from_alu(27) => 
                           write_back_op2_27_port, data_from_alu(26) => 
                           write_back_op2_26_port, data_from_alu(25) => 
                           write_back_op2_25_port, data_from_alu(24) => 
                           write_back_op2_24_port, data_from_alu(23) => 
                           write_back_op2_23_port, data_from_alu(22) => 
                           write_back_op2_22_port, data_from_alu(21) => 
                           write_back_op2_21_port, data_from_alu(20) => 
                           write_back_op2_20_port, data_from_alu(19) => 
                           write_back_op2_19_port, data_from_alu(18) => 
                           write_back_op2_18_port, data_from_alu(17) => 
                           write_back_op2_17_port, data_from_alu(16) => 
                           write_back_op2_16_port, data_from_alu(15) => 
                           write_back_op2_15_port, data_from_alu(14) => 
                           write_back_op2_14_port, data_from_alu(13) => 
                           write_back_op2_13_port, data_from_alu(12) => 
                           write_back_op2_12_port, data_from_alu(11) => 
                           write_back_op2_11_port, data_from_alu(10) => 
                           write_back_op2_10_port, data_from_alu(9) => 
                           write_back_op2_9_port, data_from_alu(8) => 
                           write_back_op2_8_port, data_from_alu(7) => 
                           write_back_op2_7_port, data_from_alu(6) => 
                           write_back_op2_6_port, data_from_alu(5) => 
                           write_back_op2_5_port, data_from_alu(4) => 
                           write_back_op2_4_port, data_from_alu(3) => 
                           write_back_op2_3_port, data_from_alu(2) => 
                           write_back_op2_2_port, data_from_alu(1) => 
                           write_back_op2_1_port, data_from_alu(0) => 
                           write_back_op2_0_port, write_back_value(31) => 
                           forward_mem_31_port, write_back_value(30) => 
                           forward_mem_30_port, write_back_value(29) => 
                           forward_mem_29_port, write_back_value(28) => 
                           forward_mem_28_port, write_back_value(27) => 
                           forward_mem_27_port, write_back_value(26) => 
                           forward_mem_26_port, write_back_value(25) => 
                           forward_mem_25_port, write_back_value(24) => 
                           forward_mem_24_port, write_back_value(23) => 
                           forward_mem_23_port, write_back_value(22) => 
                           forward_mem_22_port, write_back_value(21) => 
                           forward_mem_21_port, write_back_value(20) => 
                           forward_mem_20_port, write_back_value(19) => 
                           forward_mem_19_port, write_back_value(18) => 
                           forward_mem_18_port, write_back_value(17) => 
                           forward_mem_17_port, write_back_value(16) => 
                           forward_mem_16_port, write_back_value(15) => 
                           forward_mem_15_port, write_back_value(14) => 
                           forward_mem_14_port, write_back_value(13) => 
                           forward_mem_13_port, write_back_value(12) => 
                           forward_mem_12_port, write_back_value(11) => 
                           forward_mem_11_port, write_back_value(10) => 
                           forward_mem_10_port, write_back_value(9) => 
                           forward_mem_9_port, write_back_value(8) => 
                           forward_mem_8_port, write_back_value(7) => 
                           forward_mem_7_port, write_back_value(6) => 
                           forward_mem_6_port, write_back_value(5) => 
                           forward_mem_5_port, write_back_value(4) => 
                           forward_mem_4_port, write_back_value(3) => 
                           forward_mem_3_port, write_back_value(2) => 
                           forward_mem_2_port, write_back_value(1) => 
                           forward_mem_1_port, write_back_value(0) => 
                           forward_mem_0_port, debug(31) => debug(31), 
                           debug(30) => debug(30), debug(29) => debug(29), 
                           debug(28) => debug(28), debug(27) => debug(27), 
                           debug(26) => debug(26), debug(25) => debug(25), 
                           debug(24) => debug(24), debug(23) => debug(23), 
                           debug(22) => debug(22), debug(21) => debug(21), 
                           debug(20) => debug(20), debug(19) => debug(19), 
                           debug(18) => debug(18), debug(17) => debug(17), 
                           debug(16) => debug(16), debug(15) => debug(15), 
                           debug(14) => debug(14), debug(13) => debug(13), 
                           debug(12) => debug(12), debug(11) => debug(11), 
                           debug(10) => debug(10), debug(9) => debug(9), 
                           debug(8) => debug(8), debug(7) => debug(7), debug(6)
                           => debug(6), debug(5) => debug(5), debug(4) => 
                           debug(4), debug(3) => debug(3), debug(2) => debug(2)
                           , debug(1) => debug(1), debug(0) => debug(0));
   MU : memoryUnit port map( clock => clock, reset => reset, enable => en6, 
                           alu_result(31) => operand_res_alu_31_port, 
                           alu_result(30) => operand_res_alu_30_port, 
                           alu_result(29) => operand_res_alu_29_port, 
                           alu_result(28) => operand_res_alu_28_port, 
                           alu_result(27) => operand_res_alu_27_port, 
                           alu_result(26) => operand_res_alu_26_port, 
                           alu_result(25) => operand_res_alu_25_port, 
                           alu_result(24) => operand_res_alu_24_port, 
                           alu_result(23) => operand_res_alu_23_port, 
                           alu_result(22) => operand_res_alu_22_port, 
                           alu_result(21) => operand_res_alu_21_port, 
                           alu_result(20) => operand_res_alu_20_port, 
                           alu_result(19) => operand_res_alu_19_port, 
                           alu_result(18) => operand_res_alu_18_port, 
                           alu_result(17) => operand_res_alu_17_port, 
                           alu_result(16) => operand_res_alu_16_port, 
                           alu_result(15) => operand_res_alu_15_port, 
                           alu_result(14) => operand_res_alu_14_port, 
                           alu_result(13) => operand_res_alu_13_port, 
                           alu_result(12) => operand_res_alu_12_port, 
                           alu_result(11) => operand_res_alu_11_port, 
                           alu_result(10) => operand_res_alu_10_port, 
                           alu_result(9) => operand_res_alu_9_port, 
                           alu_result(8) => operand_res_alu_8_port, 
                           alu_result(7) => operand_res_alu_7_port, 
                           alu_result(6) => operand_res_alu_6_port, 
                           alu_result(5) => operand_res_alu_5_port, 
                           alu_result(4) => operand_res_alu_4_port, 
                           alu_result(3) => operand_res_alu_3_port, 
                           alu_result(2) => operand_res_alu_2_port, 
                           alu_result(1) => operand_res_alu_1_port, 
                           alu_result(0) => operand_res_alu_0_port, 
                           data_from_memory(31) => datain(31), 
                           data_from_memory(30) => datain(30), 
                           data_from_memory(29) => datain(29), 
                           data_from_memory(28) => datain(28), 
                           data_from_memory(27) => datain(27), 
                           data_from_memory(26) => datain(26), 
                           data_from_memory(25) => datain(25), 
                           data_from_memory(24) => datain(24), 
                           data_from_memory(23) => datain(23), 
                           data_from_memory(22) => datain(22), 
                           data_from_memory(21) => datain(21), 
                           data_from_memory(20) => datain(20), 
                           data_from_memory(19) => datain(19), 
                           data_from_memory(18) => datain(18), 
                           data_from_memory(17) => datain(17), 
                           data_from_memory(16) => datain(16), 
                           data_from_memory(15) => datain(15), 
                           data_from_memory(14) => datain(14), 
                           data_from_memory(13) => datain(13), 
                           data_from_memory(12) => datain(12), 
                           data_from_memory(11) => datain(11), 
                           data_from_memory(10) => datain(10), 
                           data_from_memory(9) => datain(9), 
                           data_from_memory(8) => datain(8), 
                           data_from_memory(7) => datain(7), 
                           data_from_memory(6) => datain(6), 
                           data_from_memory(5) => datain(5), 
                           data_from_memory(4) => datain(4), 
                           data_from_memory(3) => datain(3), 
                           data_from_memory(2) => datain(2), 
                           data_from_memory(1) => datain(1), 
                           data_from_memory(0) => datain(0), EX_MEM_Rd(4) => 
                           EX_MEM_RD_4_port, EX_MEM_Rd(3) => EX_MEM_RD_3_port, 
                           EX_MEM_Rd(2) => EX_MEM_RD_2_port, EX_MEM_Rd(1) => 
                           EX_MEM_RD_1_port, EX_MEM_Rd(0) => EX_MEM_RD_0_port, 
                           address_memory(31) => address_data_memory(31), 
                           address_memory(30) => address_data_memory(30), 
                           address_memory(29) => address_data_memory(29), 
                           address_memory(28) => address_data_memory(28), 
                           address_memory(27) => address_data_memory(27), 
                           address_memory(26) => address_data_memory(26), 
                           address_memory(25) => address_data_memory(25), 
                           address_memory(24) => address_data_memory(24), 
                           address_memory(23) => address_data_memory(23), 
                           address_memory(22) => address_data_memory(22), 
                           address_memory(21) => address_data_memory(21), 
                           address_memory(20) => address_data_memory(20), 
                           address_memory(19) => address_data_memory(19), 
                           address_memory(18) => address_data_memory(18), 
                           address_memory(17) => address_data_memory(17), 
                           address_memory(16) => address_data_memory(16), 
                           address_memory(15) => address_data_memory(15), 
                           address_memory(14) => address_data_memory(14), 
                           address_memory(13) => address_data_memory(13), 
                           address_memory(12) => address_data_memory(12), 
                           address_memory(11) => address_data_memory(11), 
                           address_memory(10) => address_data_memory(10), 
                           address_memory(9) => address_data_memory(9), 
                           address_memory(8) => address_data_memory(8), 
                           address_memory(7) => address_data_memory(7), 
                           address_memory(6) => address_data_memory(6), 
                           address_memory(5) => address_data_memory(5), 
                           address_memory(4) => address_data_memory(4), 
                           address_memory(3) => address_data_memory(3), 
                           address_memory(2) => address_data_memory(2), 
                           address_memory(1) => address_data_memory(1), 
                           address_memory(0) => address_data_memory(0), 
                           data_op1(31) => write_back_op1_31_port, data_op1(30)
                           => write_back_op1_30_port, data_op1(29) => 
                           write_back_op1_29_port, data_op1(28) => 
                           write_back_op1_28_port, data_op1(27) => 
                           write_back_op1_27_port, data_op1(26) => 
                           write_back_op1_26_port, data_op1(25) => 
                           write_back_op1_25_port, data_op1(24) => 
                           write_back_op1_24_port, data_op1(23) => 
                           write_back_op1_23_port, data_op1(22) => 
                           write_back_op1_22_port, data_op1(21) => 
                           write_back_op1_21_port, data_op1(20) => 
                           write_back_op1_20_port, data_op1(19) => 
                           write_back_op1_19_port, data_op1(18) => 
                           write_back_op1_18_port, data_op1(17) => 
                           write_back_op1_17_port, data_op1(16) => 
                           write_back_op1_16_port, data_op1(15) => 
                           write_back_op1_15_port, data_op1(14) => 
                           write_back_op1_14_port, data_op1(13) => 
                           write_back_op1_13_port, data_op1(12) => 
                           write_back_op1_12_port, data_op1(11) => 
                           write_back_op1_11_port, data_op1(10) => 
                           write_back_op1_10_port, data_op1(9) => 
                           write_back_op1_9_port, data_op1(8) => 
                           write_back_op1_8_port, data_op1(7) => 
                           write_back_op1_7_port, data_op1(6) => 
                           write_back_op1_6_port, data_op1(5) => 
                           write_back_op1_5_port, data_op1(4) => 
                           write_back_op1_4_port, data_op1(3) => 
                           write_back_op1_3_port, data_op1(2) => 
                           write_back_op1_2_port, data_op1(1) => 
                           write_back_op1_1_port, data_op1(0) => 
                           write_back_op1_0_port, data_op2(31) => 
                           write_back_op2_31_port, data_op2(30) => 
                           write_back_op2_30_port, data_op2(29) => 
                           write_back_op2_29_port, data_op2(28) => 
                           write_back_op2_28_port, data_op2(27) => 
                           write_back_op2_27_port, data_op2(26) => 
                           write_back_op2_26_port, data_op2(25) => 
                           write_back_op2_25_port, data_op2(24) => 
                           write_back_op2_24_port, data_op2(23) => 
                           write_back_op2_23_port, data_op2(22) => 
                           write_back_op2_22_port, data_op2(21) => 
                           write_back_op2_21_port, data_op2(20) => 
                           write_back_op2_20_port, data_op2(19) => 
                           write_back_op2_19_port, data_op2(18) => 
                           write_back_op2_18_port, data_op2(17) => 
                           write_back_op2_17_port, data_op2(16) => 
                           write_back_op2_16_port, data_op2(15) => 
                           write_back_op2_15_port, data_op2(14) => 
                           write_back_op2_14_port, data_op2(13) => 
                           write_back_op2_13_port, data_op2(12) => 
                           write_back_op2_12_port, data_op2(11) => 
                           write_back_op2_11_port, data_op2(10) => 
                           write_back_op2_10_port, data_op2(9) => 
                           write_back_op2_9_port, data_op2(8) => 
                           write_back_op2_8_port, data_op2(7) => 
                           write_back_op2_7_port, data_op2(6) => 
                           write_back_op2_6_port, data_op2(5) => 
                           write_back_op2_5_port, data_op2(4) => 
                           write_back_op2_4_port, data_op2(3) => 
                           write_back_op2_3_port, data_op2(2) => 
                           write_back_op2_2_port, data_op2(1) => 
                           write_back_op2_1_port, data_op2(0) => 
                           write_back_op2_0_port, MEM_WB_Rd(4) => 
                           MEM_WB_RD_4_port, MEM_WB_Rd(3) => MEM_WB_RD_3_port, 
                           MEM_WB_Rd(2) => MEM_WB_RD_2_port, MEM_WB_Rd(1) => 
                           MEM_WB_RD_1_port, MEM_WB_Rd(0) => MEM_WB_RD_0_port);
   EU : executionUnit port map( clock => clock, reset => reset, operand_a(31) 
                           => operand_A_31_port, operand_a(30) => 
                           operand_A_30_port, operand_a(29) => 
                           operand_A_29_port, operand_a(28) => 
                           operand_A_28_port, operand_a(27) => 
                           operand_A_27_port, operand_a(26) => 
                           operand_A_26_port, operand_a(25) => 
                           operand_A_25_port, operand_a(24) => 
                           operand_A_24_port, operand_a(23) => 
                           operand_A_23_port, operand_a(22) => 
                           operand_A_22_port, operand_a(21) => 
                           operand_A_21_port, operand_a(20) => 
                           operand_A_20_port, operand_a(19) => 
                           operand_A_19_port, operand_a(18) => 
                           operand_A_18_port, operand_a(17) => 
                           operand_A_17_port, operand_a(16) => 
                           operand_A_16_port, operand_a(15) => 
                           operand_A_15_port, operand_a(14) => 
                           operand_A_14_port, operand_a(13) => 
                           operand_A_13_port, operand_a(12) => 
                           operand_A_12_port, operand_a(11) => 
                           operand_A_11_port, operand_a(10) => 
                           operand_A_10_port, operand_a(9) => operand_A_9_port,
                           operand_a(8) => operand_A_8_port, operand_a(7) => 
                           operand_A_7_port, operand_a(6) => operand_A_6_port, 
                           operand_a(5) => operand_A_5_port, operand_a(4) => 
                           operand_A_4_port, operand_a(3) => operand_A_3_port, 
                           operand_a(2) => operand_A_2_port, operand_a(1) => 
                           operand_A_1_port, operand_a(0) => operand_A_0_port, 
                           operand_b(31) => operand_B_31_port, operand_b(30) =>
                           operand_B_30_port, operand_b(29) => 
                           operand_B_29_port, operand_b(28) => 
                           operand_B_28_port, operand_b(27) => 
                           operand_B_27_port, operand_b(26) => 
                           operand_B_26_port, operand_b(25) => 
                           operand_B_25_port, operand_b(24) => 
                           operand_B_24_port, operand_b(23) => 
                           operand_B_23_port, operand_b(22) => 
                           operand_B_22_port, operand_b(21) => 
                           operand_B_21_port, operand_b(20) => 
                           operand_B_20_port, operand_b(19) => 
                           operand_B_19_port, operand_b(18) => 
                           operand_B_18_port, operand_b(17) => 
                           operand_B_17_port, operand_b(16) => 
                           operand_B_16_port, operand_b(15) => 
                           operand_B_15_port, operand_b(14) => 
                           operand_B_14_port, operand_b(13) => 
                           operand_B_13_port, operand_b(12) => 
                           operand_B_12_port, operand_b(11) => 
                           operand_B_11_port, operand_b(10) => 
                           operand_B_10_port, operand_b(9) => operand_B_9_port,
                           operand_b(8) => operand_B_8_port, operand_b(7) => 
                           operand_B_7_port, operand_b(6) => operand_B_6_port, 
                           operand_b(5) => operand_B_5_port, operand_b(4) => 
                           operand_B_4_port, operand_b(3) => operand_B_3_port, 
                           operand_b(2) => operand_B_2_port, operand_b(1) => 
                           operand_B_1_port, operand_b(0) => operand_B_0_port, 
                           operand_imm(31) => operand_IMM_31_port, 
                           operand_imm(30) => operand_IMM_30_port, 
                           operand_imm(29) => operand_IMM_29_port, 
                           operand_imm(28) => operand_IMM_28_port, 
                           operand_imm(27) => operand_IMM_27_port, 
                           operand_imm(26) => operand_IMM_26_port, 
                           operand_imm(25) => operand_IMM_25_port, 
                           operand_imm(24) => operand_IMM_24_port, 
                           operand_imm(23) => operand_IMM_23_port, 
                           operand_imm(22) => operand_IMM_22_port, 
                           operand_imm(21) => operand_IMM_21_port, 
                           operand_imm(20) => operand_IMM_20_port, 
                           operand_imm(19) => operand_IMM_19_port, 
                           operand_imm(18) => operand_IMM_18_port, 
                           operand_imm(17) => operand_IMM_17_port, 
                           operand_imm(16) => operand_IMM_16_port, 
                           operand_imm(15) => operand_IMM_15_port, 
                           operand_imm(14) => operand_IMM_14_port, 
                           operand_imm(13) => operand_IMM_13_port, 
                           operand_imm(12) => operand_IMM_12_port, 
                           operand_imm(11) => operand_IMM_11_port, 
                           operand_imm(10) => operand_IMM_10_port, 
                           operand_imm(9) => operand_IMM_9_port, operand_imm(8)
                           => operand_IMM_8_port, operand_imm(7) => 
                           operand_IMM_7_port, operand_imm(6) => 
                           operand_IMM_6_port, operand_imm(5) => 
                           operand_IMM_5_port, operand_imm(4) => 
                           operand_IMM_4_port, operand_imm(3) => 
                           operand_IMM_3_port, operand_imm(2) => 
                           operand_IMM_2_port, operand_imm(1) => 
                           operand_IMM_1_port, operand_imm(0) => 
                           operand_IMM_0_port, operand_pc(31) => 
                           operand_PC_31_port, operand_pc(30) => 
                           operand_PC_30_port, operand_pc(29) => 
                           operand_PC_29_port, operand_pc(28) => 
                           operand_PC_28_port, operand_pc(27) => 
                           operand_PC_27_port, operand_pc(26) => 
                           operand_PC_26_port, operand_pc(25) => 
                           operand_PC_25_port, operand_pc(24) => 
                           operand_PC_24_port, operand_pc(23) => 
                           operand_PC_23_port, operand_pc(22) => 
                           operand_PC_22_port, operand_pc(21) => 
                           operand_PC_21_port, operand_pc(20) => 
                           operand_PC_20_port, operand_pc(19) => 
                           operand_PC_19_port, operand_pc(18) => 
                           operand_PC_18_port, operand_pc(17) => 
                           operand_PC_17_port, operand_pc(16) => 
                           operand_PC_16_port, operand_pc(15) => 
                           operand_PC_15_port, operand_pc(14) => 
                           operand_PC_14_port, operand_pc(13) => 
                           operand_PC_13_port, operand_pc(12) => 
                           operand_PC_12_port, operand_pc(11) => 
                           operand_PC_11_port, operand_pc(10) => 
                           operand_PC_10_port, operand_pc(9) => 
                           operand_PC_9_port, operand_pc(8) => 
                           operand_PC_8_port, operand_pc(7) => 
                           operand_PC_7_port, operand_pc(6) => 
                           operand_PC_6_port, operand_pc(5) => 
                           operand_PC_5_port, operand_pc(4) => 
                           operand_PC_4_port, operand_pc(3) => 
                           operand_PC_3_port, operand_pc(2) => 
                           operand_PC_2_port, operand_pc(1) => 
                           operand_PC_1_port, operand_pc(0) => 
                           operand_PC_0_port, forward_exe(31) => 
                           operand_res_alu_31_port, forward_exe(30) => 
                           operand_res_alu_30_port, forward_exe(29) => 
                           operand_res_alu_29_port, forward_exe(28) => 
                           operand_res_alu_28_port, forward_exe(27) => 
                           operand_res_alu_27_port, forward_exe(26) => 
                           operand_res_alu_26_port, forward_exe(25) => 
                           operand_res_alu_25_port, forward_exe(24) => 
                           operand_res_alu_24_port, forward_exe(23) => 
                           operand_res_alu_23_port, forward_exe(22) => 
                           operand_res_alu_22_port, forward_exe(21) => 
                           operand_res_alu_21_port, forward_exe(20) => 
                           operand_res_alu_20_port, forward_exe(19) => 
                           operand_res_alu_19_port, forward_exe(18) => 
                           operand_res_alu_18_port, forward_exe(17) => 
                           operand_res_alu_17_port, forward_exe(16) => 
                           operand_res_alu_16_port, forward_exe(15) => 
                           operand_res_alu_15_port, forward_exe(14) => 
                           operand_res_alu_14_port, forward_exe(13) => 
                           operand_res_alu_13_port, forward_exe(12) => 
                           operand_res_alu_12_port, forward_exe(11) => 
                           operand_res_alu_11_port, forward_exe(10) => 
                           operand_res_alu_10_port, forward_exe(9) => 
                           operand_res_alu_9_port, forward_exe(8) => 
                           operand_res_alu_8_port, forward_exe(7) => 
                           operand_res_alu_7_port, forward_exe(6) => 
                           operand_res_alu_6_port, forward_exe(5) => 
                           operand_res_alu_5_port, forward_exe(4) => 
                           operand_res_alu_4_port, forward_exe(3) => 
                           operand_res_alu_3_port, forward_exe(2) => 
                           operand_res_alu_2_port, forward_exe(1) => 
                           operand_res_alu_1_port, forward_exe(0) => 
                           operand_res_alu_0_port, forward_mem(31) => 
                           forward_mem_31_port, forward_mem(30) => 
                           forward_mem_30_port, forward_mem(29) => 
                           forward_mem_29_port, forward_mem(28) => 
                           forward_mem_28_port, forward_mem(27) => 
                           forward_mem_27_port, forward_mem(26) => 
                           forward_mem_26_port, forward_mem(25) => 
                           forward_mem_25_port, forward_mem(24) => 
                           forward_mem_24_port, forward_mem(23) => 
                           forward_mem_23_port, forward_mem(22) => 
                           forward_mem_22_port, forward_mem(21) => 
                           forward_mem_21_port, forward_mem(20) => 
                           forward_mem_20_port, forward_mem(19) => 
                           forward_mem_19_port, forward_mem(18) => 
                           forward_mem_18_port, forward_mem(17) => 
                           forward_mem_17_port, forward_mem(16) => 
                           forward_mem_16_port, forward_mem(15) => 
                           forward_mem_15_port, forward_mem(14) => 
                           forward_mem_14_port, forward_mem(13) => 
                           forward_mem_13_port, forward_mem(12) => 
                           forward_mem_12_port, forward_mem(11) => 
                           forward_mem_11_port, forward_mem(10) => 
                           forward_mem_10_port, forward_mem(9) => 
                           forward_mem_9_port, forward_mem(8) => 
                           forward_mem_8_port, forward_mem(7) => 
                           forward_mem_7_port, forward_mem(6) => 
                           forward_mem_6_port, forward_mem(5) => 
                           forward_mem_5_port, forward_mem(4) => 
                           forward_mem_4_port, forward_mem(3) => 
                           forward_mem_3_port, forward_mem(2) => 
                           forward_mem_2_port, forward_mem(1) => 
                           forward_mem_1_port, forward_mem(0) => 
                           forward_mem_0_port, EX_MEM_write => EX_MEM_write, 
                           MEM_WB_write => MEM_WB_write, MEM_WB_rd(4) => 
                           MEM_WB_RD_4_port, MEM_WB_rd(3) => MEM_WB_RD_3_port, 
                           MEM_WB_rd(2) => MEM_WB_RD_2_port, MEM_WB_rd(1) => 
                           MEM_WB_RD_1_port, MEM_WB_rd(0) => MEM_WB_RD_0_port, 
                           ID_EX_Rd(4) => ID_EX_Rd_4_port, ID_EX_Rd(3) => 
                           ID_EX_Rd_3_port, ID_EX_Rd(2) => ID_EX_Rd_2_port, 
                           ID_EX_Rd(1) => ID_EX_Rd_1_port, ID_EX_Rd(0) => 
                           ID_EX_Rd_0_port, ID_EX_Rs(4) => ID_EX_Rs_4_port, 
                           ID_EX_Rs(3) => ID_EX_Rs_3_port, ID_EX_Rs(2) => 
                           ID_EX_Rs_2_port, ID_EX_Rs(1) => ID_EX_Rs_1_port, 
                           ID_EX_Rs(0) => ID_EX_Rs_0_port, ID_EX_Rt(4) => 
                           ID_EX_Rt_4_port, ID_EX_Rt(3) => ID_EX_Rt_3_port, 
                           ID_EX_Rt(2) => ID_EX_Rt_2_port, ID_EX_Rt(1) => 
                           ID_EX_Rt_1_port, ID_EX_Rt(0) => ID_EX_Rt_0_port, 
                           enable => en5, sel_1 => sel1, sel_2 => sel2, sel_3 
                           => sel3, func(10) => func(10), func(9) => func(9), 
                           func(8) => func(8), func(7) => func(7), func(6) => 
                           func(6), func(5) => func(5), func(4) => func(4), 
                           func(3) => func(3), func(2) => func(2), func(1) => 
                           func(1), func(0) => func(0), EX_MEM_rd(4) => 
                           EX_MEM_RD_4_port, EX_MEM_rd(3) => EX_MEM_RD_3_port, 
                           EX_MEM_rd(2) => EX_MEM_RD_2_port, EX_MEM_rd(1) => 
                           EX_MEM_RD_1_port, EX_MEM_rd(0) => EX_MEM_RD_0_port, 
                           out_res_operand_one(31) => operand_res_alu_31_port, 
                           out_res_operand_one(30) => operand_res_alu_30_port, 
                           out_res_operand_one(29) => operand_res_alu_29_port, 
                           out_res_operand_one(28) => operand_res_alu_28_port, 
                           out_res_operand_one(27) => operand_res_alu_27_port, 
                           out_res_operand_one(26) => operand_res_alu_26_port, 
                           out_res_operand_one(25) => operand_res_alu_25_port, 
                           out_res_operand_one(24) => operand_res_alu_24_port, 
                           out_res_operand_one(23) => operand_res_alu_23_port, 
                           out_res_operand_one(22) => operand_res_alu_22_port, 
                           out_res_operand_one(21) => operand_res_alu_21_port, 
                           out_res_operand_one(20) => operand_res_alu_20_port, 
                           out_res_operand_one(19) => operand_res_alu_19_port, 
                           out_res_operand_one(18) => operand_res_alu_18_port, 
                           out_res_operand_one(17) => operand_res_alu_17_port, 
                           out_res_operand_one(16) => operand_res_alu_16_port, 
                           out_res_operand_one(15) => operand_res_alu_15_port, 
                           out_res_operand_one(14) => operand_res_alu_14_port, 
                           out_res_operand_one(13) => operand_res_alu_13_port, 
                           out_res_operand_one(12) => operand_res_alu_12_port, 
                           out_res_operand_one(11) => operand_res_alu_11_port, 
                           out_res_operand_one(10) => operand_res_alu_10_port, 
                           out_res_operand_one(9) => operand_res_alu_9_port, 
                           out_res_operand_one(8) => operand_res_alu_8_port, 
                           out_res_operand_one(7) => operand_res_alu_7_port, 
                           out_res_operand_one(6) => operand_res_alu_6_port, 
                           out_res_operand_one(5) => operand_res_alu_5_port, 
                           out_res_operand_one(4) => operand_res_alu_4_port, 
                           out_res_operand_one(3) => operand_res_alu_3_port, 
                           out_res_operand_one(2) => operand_res_alu_2_port, 
                           out_res_operand_one(1) => operand_res_alu_1_port, 
                           out_res_operand_one(0) => operand_res_alu_0_port, 
                           out_res_operand_two(31) => dataout(31), 
                           out_res_operand_two(30) => dataout(30), 
                           out_res_operand_two(29) => dataout(29), 
                           out_res_operand_two(28) => dataout(28), 
                           out_res_operand_two(27) => dataout(27), 
                           out_res_operand_two(26) => dataout(26), 
                           out_res_operand_two(25) => dataout(25), 
                           out_res_operand_two(24) => dataout(24), 
                           out_res_operand_two(23) => dataout(23), 
                           out_res_operand_two(22) => dataout(22), 
                           out_res_operand_two(21) => dataout(21), 
                           out_res_operand_two(20) => dataout(20), 
                           out_res_operand_two(19) => dataout(19), 
                           out_res_operand_two(18) => dataout(18), 
                           out_res_operand_two(17) => dataout(17), 
                           out_res_operand_two(16) => dataout(16), 
                           out_res_operand_two(15) => dataout(15), 
                           out_res_operand_two(14) => dataout(14), 
                           out_res_operand_two(13) => dataout(13), 
                           out_res_operand_two(12) => dataout(12), 
                           out_res_operand_two(11) => dataout(11), 
                           out_res_operand_two(10) => dataout(10), 
                           out_res_operand_two(9) => dataout(9), 
                           out_res_operand_two(8) => dataout(8), 
                           out_res_operand_two(7) => dataout(7), 
                           out_res_operand_two(6) => dataout(6), 
                           out_res_operand_two(5) => dataout(5), 
                           out_res_operand_two(4) => dataout(4), 
                           out_res_operand_two(3) => dataout(3), 
                           out_res_operand_two(2) => dataout(2), 
                           out_res_operand_two(1) => dataout(1), 
                           out_res_operand_two(0) => dataout(0), next_pc(31) =>
                           next_pc_31_port, next_pc(30) => next_pc_30_port, 
                           next_pc(29) => next_pc_29_port, next_pc(28) => 
                           next_pc_28_port, next_pc(27) => next_pc_27_port, 
                           next_pc(26) => next_pc_26_port, next_pc(25) => 
                           next_pc_25_port, next_pc(24) => next_pc_24_port, 
                           next_pc(23) => next_pc_23_port, next_pc(22) => 
                           next_pc_22_port, next_pc(21) => next_pc_21_port, 
                           next_pc(20) => next_pc_20_port, next_pc(19) => 
                           next_pc_19_port, next_pc(18) => next_pc_18_port, 
                           next_pc(17) => next_pc_17_port, next_pc(16) => 
                           next_pc_16_port, next_pc(15) => next_pc_15_port, 
                           next_pc(14) => next_pc_14_port, next_pc(13) => 
                           next_pc_13_port, next_pc(12) => next_pc_12_port, 
                           next_pc(11) => next_pc_11_port, next_pc(10) => 
                           next_pc_10_port, next_pc(9) => next_pc_9_port, 
                           next_pc(8) => next_pc_8_port, next_pc(7) => 
                           next_pc_7_port, next_pc(6) => next_pc_6_port, 
                           next_pc(5) => next_pc_5_port, next_pc(4) => 
                           next_pc_4_port, next_pc(3) => next_pc_3_port, 
                           next_pc(2) => next_pc_2_port, next_pc(1) => 
                           next_pc_1_port, next_pc(0) => next_pc_0_port, jump 
                           => jump, multi_cycle_operation => 
                           multi_cycle_operation);
   DU : decodeUnit port map( clock => clock, reset => reset, en1 => en1, 
                           read_enable_portA => en2, read_enable_portB => en3, 
                           write_enable_portW => en4, instructionWord(31) => 
                           instruction_31_port, instructionWord(30) => 
                           instruction_30_port, instructionWord(29) => 
                           instruction_29_port, instructionWord(28) => 
                           instruction_28_port, instructionWord(27) => 
                           instruction_27_port, instructionWord(26) => 
                           instruction_26_port, instructionWord(25) => 
                           instruction_25_port, instructionWord(24) => 
                           instruction_24_port, instructionWord(23) => 
                           instruction_23_port, instructionWord(22) => 
                           instruction_22_port, instructionWord(21) => 
                           instruction_21_port, instructionWord(20) => 
                           instruction_20_port, instructionWord(19) => 
                           instruction_19_port, instructionWord(18) => 
                           instruction_18_port, instructionWord(17) => 
                           instruction_17_port, instructionWord(16) => 
                           instruction_16_port, instructionWord(15) => 
                           instruction_15_port, instructionWord(14) => 
                           instruction_14_port, instructionWord(13) => 
                           instruction_13_port, instructionWord(12) => 
                           instruction_12_port, instructionWord(11) => 
                           instruction_11_port, instructionWord(10) => 
                           instruction_10_port, instructionWord(9) => 
                           instruction_9_port, instructionWord(8) => 
                           instruction_8_port, instructionWord(7) => 
                           instruction_7_port, instructionWord(6) => 
                           instruction_6_port, instructionWord(5) => 
                           instruction_5_port, instructionWord(4) => 
                           instruction_4_port, instructionWord(3) => 
                           instruction_3_port, instructionWord(2) => 
                           instruction_2_port, instructionWord(1) => 
                           instruction_1_port, instructionWord(0) => 
                           instruction_0_port, ID_EX_MemRead => 
                           hazard_condition, ID_EX_RT_Address(4) => 
                           ID_EX_Rt_4_port, ID_EX_RT_Address(3) => 
                           ID_EX_Rt_3_port, ID_EX_RT_Address(2) => 
                           ID_EX_Rt_2_port, ID_EX_RT_Address(1) => 
                           ID_EX_Rt_1_port, ID_EX_RT_Address(0) => 
                           ID_EX_Rt_0_port, writeData(31) => 
                           forward_mem_31_port, writeData(30) => 
                           forward_mem_30_port, writeData(29) => 
                           forward_mem_29_port, writeData(28) => 
                           forward_mem_28_port, writeData(27) => 
                           forward_mem_27_port, writeData(26) => 
                           forward_mem_26_port, writeData(25) => 
                           forward_mem_25_port, writeData(24) => 
                           forward_mem_24_port, writeData(23) => 
                           forward_mem_23_port, writeData(22) => 
                           forward_mem_22_port, writeData(21) => 
                           forward_mem_21_port, writeData(20) => 
                           forward_mem_20_port, writeData(19) => 
                           forward_mem_19_port, writeData(18) => 
                           forward_mem_18_port, writeData(17) => 
                           forward_mem_17_port, writeData(16) => 
                           forward_mem_16_port, writeData(15) => 
                           forward_mem_15_port, writeData(14) => 
                           forward_mem_14_port, writeData(13) => 
                           forward_mem_13_port, writeData(12) => 
                           forward_mem_12_port, writeData(11) => 
                           forward_mem_11_port, writeData(10) => 
                           forward_mem_10_port, writeData(9) => 
                           forward_mem_9_port, writeData(8) => 
                           forward_mem_8_port, writeData(7) => 
                           forward_mem_7_port, writeData(6) => 
                           forward_mem_6_port, writeData(5) => 
                           forward_mem_5_port, writeData(4) => 
                           forward_mem_4_port, writeData(3) => 
                           forward_mem_3_port, writeData(2) => 
                           forward_mem_2_port, writeData(1) => 
                           forward_mem_1_port, writeData(0) => 
                           forward_mem_0_port, writeAddress(4) => 
                           MEM_WB_RD_4_port, writeAddress(3) => 
                           MEM_WB_RD_3_port, writeAddress(2) => 
                           MEM_WB_RD_2_port, writeAddress(1) => 
                           MEM_WB_RD_1_port, writeAddress(0) => 
                           MEM_WB_RD_0_port, pc(31) => NPC_to_decode_31_port, 
                           pc(30) => NPC_to_decode_30_port, pc(29) => 
                           NPC_to_decode_29_port, pc(28) => 
                           NPC_to_decode_28_port, pc(27) => 
                           NPC_to_decode_27_port, pc(26) => 
                           NPC_to_decode_26_port, pc(25) => 
                           NPC_to_decode_25_port, pc(24) => 
                           NPC_to_decode_24_port, pc(23) => 
                           NPC_to_decode_23_port, pc(22) => 
                           NPC_to_decode_22_port, pc(21) => 
                           NPC_to_decode_21_port, pc(20) => 
                           NPC_to_decode_20_port, pc(19) => 
                           NPC_to_decode_19_port, pc(18) => 
                           NPC_to_decode_18_port, pc(17) => 
                           NPC_to_decode_17_port, pc(16) => 
                           NPC_to_decode_16_port, pc(15) => 
                           NPC_to_decode_15_port, pc(14) => 
                           NPC_to_decode_14_port, pc(13) => 
                           NPC_to_decode_13_port, pc(12) => 
                           NPC_to_decode_12_port, pc(11) => 
                           NPC_to_decode_11_port, pc(10) => 
                           NPC_to_decode_10_port, pc(9) => NPC_to_decode_9_port
                           , pc(8) => NPC_to_decode_8_port, pc(7) => 
                           NPC_to_decode_7_port, pc(6) => NPC_to_decode_6_port,
                           pc(5) => NPC_to_decode_5_port, pc(4) => 
                           NPC_to_decode_4_port, pc(3) => NPC_to_decode_3_port,
                           pc(2) => NPC_to_decode_2_port, pc(1) => 
                           NPC_to_decode_1_port, pc(0) => NPC_to_decode_0_port,
                           sel_ext => sel_ext, multi_cycle_operation => 
                           multi_cycle_operation, enable_signal_PC_IF_ID => 
                           disable_fetch_register, selectNop => hazard_detected
                           , outRT(4) => ID_EX_Rt_4_port, outRT(3) => 
                           ID_EX_Rt_3_port, outRT(2) => ID_EX_Rt_2_port, 
                           outRT(1) => ID_EX_Rt_1_port, outRT(0) => 
                           ID_EX_Rt_0_port, outRD(4) => ID_EX_Rd_4_port, 
                           outRD(3) => ID_EX_Rd_3_port, outRD(2) => 
                           ID_EX_Rd_2_port, outRD(1) => ID_EX_Rd_1_port, 
                           outRD(0) => ID_EX_Rd_0_port, outRS(4) => 
                           ID_EX_Rs_4_port, outRS(3) => ID_EX_Rs_3_port, 
                           outRS(2) => ID_EX_Rs_2_port, outRS(1) => 
                           ID_EX_Rs_1_port, outRS(0) => ID_EX_Rs_0_port, 
                           outIMM(31) => operand_IMM_31_port, outIMM(30) => 
                           operand_IMM_30_port, outIMM(29) => 
                           operand_IMM_29_port, outIMM(28) => 
                           operand_IMM_28_port, outIMM(27) => 
                           operand_IMM_27_port, outIMM(26) => 
                           operand_IMM_26_port, outIMM(25) => 
                           operand_IMM_25_port, outIMM(24) => 
                           operand_IMM_24_port, outIMM(23) => 
                           operand_IMM_23_port, outIMM(22) => 
                           operand_IMM_22_port, outIMM(21) => 
                           operand_IMM_21_port, outIMM(20) => 
                           operand_IMM_20_port, outIMM(19) => 
                           operand_IMM_19_port, outIMM(18) => 
                           operand_IMM_18_port, outIMM(17) => 
                           operand_IMM_17_port, outIMM(16) => 
                           operand_IMM_16_port, outIMM(15) => 
                           operand_IMM_15_port, outIMM(14) => 
                           operand_IMM_14_port, outIMM(13) => 
                           operand_IMM_13_port, outIMM(12) => 
                           operand_IMM_12_port, outIMM(11) => 
                           operand_IMM_11_port, outIMM(10) => 
                           operand_IMM_10_port, outIMM(9) => operand_IMM_9_port
                           , outIMM(8) => operand_IMM_8_port, outIMM(7) => 
                           operand_IMM_7_port, outIMM(6) => operand_IMM_6_port,
                           outIMM(5) => operand_IMM_5_port, outIMM(4) => 
                           operand_IMM_4_port, outIMM(3) => operand_IMM_3_port,
                           outIMM(2) => operand_IMM_2_port, outIMM(1) => 
                           operand_IMM_1_port, outIMM(0) => operand_IMM_0_port,
                           outPC(31) => operand_PC_31_port, outPC(30) => 
                           operand_PC_30_port, outPC(29) => operand_PC_29_port,
                           outPC(28) => operand_PC_28_port, outPC(27) => 
                           operand_PC_27_port, outPC(26) => operand_PC_26_port,
                           outPC(25) => operand_PC_25_port, outPC(24) => 
                           operand_PC_24_port, outPC(23) => operand_PC_23_port,
                           outPC(22) => operand_PC_22_port, outPC(21) => 
                           operand_PC_21_port, outPC(20) => operand_PC_20_port,
                           outPC(19) => operand_PC_19_port, outPC(18) => 
                           operand_PC_18_port, outPC(17) => operand_PC_17_port,
                           outPC(16) => operand_PC_16_port, outPC(15) => 
                           operand_PC_15_port, outPC(14) => operand_PC_14_port,
                           outPC(13) => operand_PC_13_port, outPC(12) => 
                           operand_PC_12_port, outPC(11) => operand_PC_11_port,
                           outPC(10) => operand_PC_10_port, outPC(9) => 
                           operand_PC_9_port, outPC(8) => operand_PC_8_port, 
                           outPC(7) => operand_PC_7_port, outPC(6) => 
                           operand_PC_6_port, outPC(5) => operand_PC_5_port, 
                           outPC(4) => operand_PC_4_port, outPC(3) => 
                           operand_PC_3_port, outPC(2) => operand_PC_2_port, 
                           outPC(1) => operand_PC_1_port, outPC(0) => 
                           operand_PC_0_port, outA(31) => operand_A_31_port, 
                           outA(30) => operand_A_30_port, outA(29) => 
                           operand_A_29_port, outA(28) => operand_A_28_port, 
                           outA(27) => operand_A_27_port, outA(26) => 
                           operand_A_26_port, outA(25) => operand_A_25_port, 
                           outA(24) => operand_A_24_port, outA(23) => 
                           operand_A_23_port, outA(22) => operand_A_22_port, 
                           outA(21) => operand_A_21_port, outA(20) => 
                           operand_A_20_port, outA(19) => operand_A_19_port, 
                           outA(18) => operand_A_18_port, outA(17) => 
                           operand_A_17_port, outA(16) => operand_A_16_port, 
                           outA(15) => operand_A_15_port, outA(14) => 
                           operand_A_14_port, outA(13) => operand_A_13_port, 
                           outA(12) => operand_A_12_port, outA(11) => 
                           operand_A_11_port, outA(10) => operand_A_10_port, 
                           outA(9) => operand_A_9_port, outA(8) => 
                           operand_A_8_port, outA(7) => operand_A_7_port, 
                           outA(6) => operand_A_6_port, outA(5) => 
                           operand_A_5_port, outA(4) => operand_A_4_port, 
                           outA(3) => operand_A_3_port, outA(2) => 
                           operand_A_2_port, outA(1) => operand_A_1_port, 
                           outA(0) => operand_A_0_port, outB(31) => 
                           operand_B_31_port, outB(30) => operand_B_30_port, 
                           outB(29) => operand_B_29_port, outB(28) => 
                           operand_B_28_port, outB(27) => operand_B_27_port, 
                           outB(26) => operand_B_26_port, outB(25) => 
                           operand_B_25_port, outB(24) => operand_B_24_port, 
                           outB(23) => operand_B_23_port, outB(22) => 
                           operand_B_22_port, outB(21) => operand_B_21_port, 
                           outB(20) => operand_B_20_port, outB(19) => 
                           operand_B_19_port, outB(18) => operand_B_18_port, 
                           outB(17) => operand_B_17_port, outB(16) => 
                           operand_B_16_port, outB(15) => operand_B_15_port, 
                           outB(14) => operand_B_14_port, outB(13) => 
                           operand_B_13_port, outB(12) => operand_B_12_port, 
                           outB(11) => operand_B_11_port, outB(10) => 
                           operand_B_10_port, outB(9) => operand_B_9_port, 
                           outB(8) => operand_B_8_port, outB(7) => 
                           operand_B_7_port, outB(6) => operand_B_6_port, 
                           outB(5) => operand_B_5_port, outB(4) => 
                           operand_B_4_port, outB(3) => operand_B_3_port, 
                           outB(2) => operand_B_2_port, outB(1) => 
                           operand_B_1_port, outB(0) => operand_B_0_port);
   FU : fetchUnit port map( sel0 => sel0, en0 => disable_fetch_register, clock 
                           => clock, reset => reset, fromInstructionMemory(31) 
                           => from_instruction_memory(31), 
                           fromInstructionMemory(30) => 
                           from_instruction_memory(30), 
                           fromInstructionMemory(29) => 
                           from_instruction_memory(29), 
                           fromInstructionMemory(28) => 
                           from_instruction_memory(28), 
                           fromInstructionMemory(27) => 
                           from_instruction_memory(27), 
                           fromInstructionMemory(26) => 
                           from_instruction_memory(26), 
                           fromInstructionMemory(25) => 
                           from_instruction_memory(25), 
                           fromInstructionMemory(24) => 
                           from_instruction_memory(24), 
                           fromInstructionMemory(23) => 
                           from_instruction_memory(23), 
                           fromInstructionMemory(22) => 
                           from_instruction_memory(22), 
                           fromInstructionMemory(21) => 
                           from_instruction_memory(21), 
                           fromInstructionMemory(20) => 
                           from_instruction_memory(20), 
                           fromInstructionMemory(19) => 
                           from_instruction_memory(19), 
                           fromInstructionMemory(18) => 
                           from_instruction_memory(18), 
                           fromInstructionMemory(17) => 
                           from_instruction_memory(17), 
                           fromInstructionMemory(16) => 
                           from_instruction_memory(16), 
                           fromInstructionMemory(15) => 
                           from_instruction_memory(15), 
                           fromInstructionMemory(14) => 
                           from_instruction_memory(14), 
                           fromInstructionMemory(13) => 
                           from_instruction_memory(13), 
                           fromInstructionMemory(12) => 
                           from_instruction_memory(12), 
                           fromInstructionMemory(11) => 
                           from_instruction_memory(11), 
                           fromInstructionMemory(10) => 
                           from_instruction_memory(10), 
                           fromInstructionMemory(9) => 
                           from_instruction_memory(9), fromInstructionMemory(8)
                           => from_instruction_memory(8), 
                           fromInstructionMemory(7) => 
                           from_instruction_memory(7), fromInstructionMemory(6)
                           => from_instruction_memory(6), 
                           fromInstructionMemory(5) => 
                           from_instruction_memory(5), fromInstructionMemory(4)
                           => from_instruction_memory(4), 
                           fromInstructionMemory(3) => 
                           from_instruction_memory(3), fromInstructionMemory(2)
                           => from_instruction_memory(2), 
                           fromInstructionMemory(1) => 
                           from_instruction_memory(1), fromInstructionMemory(0)
                           => from_instruction_memory(0), next_PC(31) => 
                           next_pc_31_port, next_PC(30) => next_pc_30_port, 
                           next_PC(29) => next_pc_29_port, next_PC(28) => 
                           next_pc_28_port, next_PC(27) => next_pc_27_port, 
                           next_PC(26) => next_pc_26_port, next_PC(25) => 
                           next_pc_25_port, next_PC(24) => next_pc_24_port, 
                           next_PC(23) => next_pc_23_port, next_PC(22) => 
                           next_pc_22_port, next_PC(21) => next_pc_21_port, 
                           next_PC(20) => next_pc_20_port, next_PC(19) => 
                           next_pc_19_port, next_PC(18) => next_pc_18_port, 
                           next_PC(17) => next_pc_17_port, next_PC(16) => 
                           next_pc_16_port, next_PC(15) => next_pc_15_port, 
                           next_PC(14) => next_pc_14_port, next_PC(13) => 
                           next_pc_13_port, next_PC(12) => next_pc_12_port, 
                           next_PC(11) => next_pc_11_port, next_PC(10) => 
                           next_pc_10_port, next_PC(9) => next_pc_9_port, 
                           next_PC(8) => next_pc_8_port, next_PC(7) => 
                           next_pc_7_port, next_PC(6) => next_pc_6_port, 
                           next_PC(5) => next_pc_5_port, next_PC(4) => 
                           next_pc_4_port, next_PC(3) => next_pc_3_port, 
                           next_PC(2) => next_pc_2_port, next_PC(1) => 
                           next_pc_1_port, next_PC(0) => next_pc_0_port, 
                           PcToInstructionMemory(31) => pc_to_im(31), 
                           PcToInstructionMemory(30) => pc_to_im(30), 
                           PcToInstructionMemory(29) => pc_to_im(29), 
                           PcToInstructionMemory(28) => pc_to_im(28), 
                           PcToInstructionMemory(27) => pc_to_im(27), 
                           PcToInstructionMemory(26) => pc_to_im(26), 
                           PcToInstructionMemory(25) => pc_to_im(25), 
                           PcToInstructionMemory(24) => pc_to_im(24), 
                           PcToInstructionMemory(23) => pc_to_im(23), 
                           PcToInstructionMemory(22) => pc_to_im(22), 
                           PcToInstructionMemory(21) => pc_to_im(21), 
                           PcToInstructionMemory(20) => pc_to_im(20), 
                           PcToInstructionMemory(19) => pc_to_im(19), 
                           PcToInstructionMemory(18) => pc_to_im(18), 
                           PcToInstructionMemory(17) => pc_to_im(17), 
                           PcToInstructionMemory(16) => pc_to_im(16), 
                           PcToInstructionMemory(15) => pc_to_im(15), 
                           PcToInstructionMemory(14) => pc_to_im(14), 
                           PcToInstructionMemory(13) => pc_to_im(13), 
                           PcToInstructionMemory(12) => pc_to_im(12), 
                           PcToInstructionMemory(11) => pc_to_im(11), 
                           PcToInstructionMemory(10) => pc_to_im(10), 
                           PcToInstructionMemory(9) => pc_to_im(9), 
                           PcToInstructionMemory(8) => pc_to_im(8), 
                           PcToInstructionMemory(7) => pc_to_im(7), 
                           PcToInstructionMemory(6) => pc_to_im(6), 
                           PcToInstructionMemory(5) => pc_to_im(5), 
                           PcToInstructionMemory(4) => pc_to_im(4), 
                           PcToInstructionMemory(3) => pc_to_im(3), 
                           PcToInstructionMemory(2) => pc_to_im(2), 
                           PcToInstructionMemory(1) => pc_to_im(1), 
                           PcToInstructionMemory(0) => pc_to_im(0), 
                           InstructionToDecode(31) => instruction_31_port, 
                           InstructionToDecode(30) => instruction_30_port, 
                           InstructionToDecode(29) => instruction_29_port, 
                           InstructionToDecode(28) => instruction_28_port, 
                           InstructionToDecode(27) => instruction_27_port, 
                           InstructionToDecode(26) => instruction_26_port, 
                           InstructionToDecode(25) => instruction_25_port, 
                           InstructionToDecode(24) => instruction_24_port, 
                           InstructionToDecode(23) => instruction_23_port, 
                           InstructionToDecode(22) => instruction_22_port, 
                           InstructionToDecode(21) => instruction_21_port, 
                           InstructionToDecode(20) => instruction_20_port, 
                           InstructionToDecode(19) => instruction_19_port, 
                           InstructionToDecode(18) => instruction_18_port, 
                           InstructionToDecode(17) => instruction_17_port, 
                           InstructionToDecode(16) => instruction_16_port, 
                           InstructionToDecode(15) => instruction_15_port, 
                           InstructionToDecode(14) => instruction_14_port, 
                           InstructionToDecode(13) => instruction_13_port, 
                           InstructionToDecode(12) => instruction_12_port, 
                           InstructionToDecode(11) => instruction_11_port, 
                           InstructionToDecode(10) => instruction_10_port, 
                           InstructionToDecode(9) => instruction_9_port, 
                           InstructionToDecode(8) => instruction_8_port, 
                           InstructionToDecode(7) => instruction_7_port, 
                           InstructionToDecode(6) => instruction_6_port, 
                           InstructionToDecode(5) => instruction_5_port, 
                           InstructionToDecode(4) => instruction_4_port, 
                           InstructionToDecode(3) => instruction_3_port, 
                           InstructionToDecode(2) => instruction_2_port, 
                           InstructionToDecode(1) => instruction_1_port, 
                           InstructionToDecode(0) => instruction_0_port, 
                           pcToDecode(31) => NPC_to_decode_31_port, 
                           pcToDecode(30) => NPC_to_decode_30_port, 
                           pcToDecode(29) => NPC_to_decode_29_port, 
                           pcToDecode(28) => NPC_to_decode_28_port, 
                           pcToDecode(27) => NPC_to_decode_27_port, 
                           pcToDecode(26) => NPC_to_decode_26_port, 
                           pcToDecode(25) => NPC_to_decode_25_port, 
                           pcToDecode(24) => NPC_to_decode_24_port, 
                           pcToDecode(23) => NPC_to_decode_23_port, 
                           pcToDecode(22) => NPC_to_decode_22_port, 
                           pcToDecode(21) => NPC_to_decode_21_port, 
                           pcToDecode(20) => NPC_to_decode_20_port, 
                           pcToDecode(19) => NPC_to_decode_19_port, 
                           pcToDecode(18) => NPC_to_decode_18_port, 
                           pcToDecode(17) => NPC_to_decode_17_port, 
                           pcToDecode(16) => NPC_to_decode_16_port, 
                           pcToDecode(15) => NPC_to_decode_15_port, 
                           pcToDecode(14) => NPC_to_decode_14_port, 
                           pcToDecode(13) => NPC_to_decode_13_port, 
                           pcToDecode(12) => NPC_to_decode_12_port, 
                           pcToDecode(11) => NPC_to_decode_11_port, 
                           pcToDecode(10) => NPC_to_decode_10_port, 
                           pcToDecode(9) => NPC_to_decode_9_port, pcToDecode(8)
                           => NPC_to_decode_8_port, pcToDecode(7) => 
                           NPC_to_decode_7_port, pcToDecode(6) => 
                           NPC_to_decode_6_port, pcToDecode(5) => 
                           NPC_to_decode_5_port, pcToDecode(4) => 
                           NPC_to_decode_4_port, pcToDecode(3) => 
                           NPC_to_decode_3_port, pcToDecode(2) => 
                           NPC_to_decode_2_port, pcToDecode(1) => 
                           NPC_to_decode_1_port, pcToDecode(0) => 
                           NPC_to_decode_0_port);

end SYN_Structural;
